// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
CL4RXZpXoDig50Rlw9Q/5Yv92c5h5YN84J7T9knCvt9WbFvDeq9Hm0f0mmo31xGXL5rtX/vernZG
nBebkS5qcrD8mBBLQak680/W3Al1B4ApJBgqUIFcfxct8/pd++Yutc1anIliqpWf5Tpk8NjtoDNG
dwLQBo5FKQhvEo3ecCQFPgRLc9MuxVWHqT3l1sYsGytQcnfSdyAqd66UQh64y7RVBb0Ont9/Z3sa
I6cNxVkZxurlpqDoV6H3o/3nrPrFkvaUkycaY51W/KtUXPJ3OOJhJw+kB28gpevHEjCN7V3jyxoI
XlsAMKfWh2/sYFmXBnSLbfNzGEwPEIrLM/PHnA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1SKAfP+nhMM12Vz7XUF2R+Fwlj6wVvcz2S6YSPFYmWMeg/Bjvpekb48M3S/vqt6hd7ZZ1HbWdcIF
eFhKUb6ZrtfLNeoWT9yKrJQHUFF0O4+7/Y6VPu9bBHey+aDsEKPewg6hXej0h4+9uSe6EOFQlU0n
ZqvW1GjX4dewNT6JhKqrQc/Qex9/+fmw+MXLw0HUcnKA9XIS9BW+Qp/kVOYhQa6BJ0DP3sPErOjl
f6ROL4Y29UIibYAPZUylX4Dkmq2WTLdGwTAwOqVypQlGhtXjO5TKHVTOLvqE8JVs5N34O3CWbTYU
CF6yoJ9ws6dWpqSegRdSA38gk92QhOBGjvdr7hvHC2/euHMLco4MpBh5faGNdOtjMKSo4Bxzsn32
1riXlBFDqMO40nCqBUMRk7HdcAg9bBg79HAwXu06YCIuUOfQvpM8Z0pKHjaYXCNTkQZDiMmzcAZE
CKO1e9g0yJIM9PCq2X2FTKWSLsHDeLQ37DY5lscQcS3x8a3VdgIIndDR5VnhkEnGQ/aMi3BxFIgR
qHk735HlndX9eX1ppwJbknkIW1urXXXHML7IY03eocwu1C2JMRDmk5fmBZDAdiaG8qDrVWlOZdUm
PTRzUMMWDpsZVxpp//jPQUq1aSp/SSuP6nS+xeywOtBvuN3zewEQdse05iL5hMr7VnlgGxr0zcch
sehvEM+nhaVPHbyi1nr2/dl+YS/6CpNvOf0YOjcNqkZm9Oyx5Hx4f8DHyeC0B7nCMxre/5+DZlIJ
+k3CsdiYVAPk1M+k7fjRHk+bUmUXlH+2AX15v2eLcKxlQX0Poarub9I3qXl3p0ljG55dK5Ur61Ez
pr74LnZ6mxhOfr0PtjeBDrkpXz0Aiw8NLL4gD4gxKLc8LCuCQYYj8KRzMvr6gNtYFZEAyZj1DjGt
fPkHHnUhtMt2ctb0yqP7oSlLTgYy1jSWWR3R8YwzRCb2h40RtJyF6AjWW1s3okouEr0u5aSRg+0J
9wQBgWGH4nQTB64M4KUEJp2iyEp8plBRu8lTs/79e62HnjD8V2lQIFEUf7qV7Tvl6xO/YS/2d7iD
dFh0vO8qV9eWsEcR6bSezVTobQ8Et3GroLyY8+fXtFZP1jliv/eYEAiGANZSQnbP8lBz5rqmNNJp
Ur36+1nn/ihHBqYShz5NMkYyn6rOp5HoG67hqKnqi7rk1A0kLVaSh2kwRZ2811YG4PQQgJPXxjYo
afHhv5LDrgn3aliiTPE3Xk+7/0KM20DHgO8YPD0UD9bdZcr9cf2tImMkhrim8czSNmxA/FagUdbR
FsngSqV4xJwlIcUt0bTKiLVu9YHzIj7yzlUMYTaoWoTdEj5PAkvVtC0byog2I9q9oMkjX38Ur3cu
NXVL7nycte5uglyCOA4ZOLGSJQS0dIbdoV+VXB4oGORegByEM1asQK2XwRmAlEe3uEf8zCmdXRm3
RjtyQhNdrry/VOG7iPAkEXFCLjw6YP9QfF2IwwmgmwS/kORiTmzNmCu1rHt3ktu2PQNxDK5kKEdM
W90IcguUhBbDCEtNJqv+ZKArA1xkabGo0mwgf8vcDNmpHh6jR8jh89yO5gLQoar0WGw2xoFlh9n0
2kygaZ6J65Flv/54zcpAy7qpZy+89blY81H82pyS6fyx+YLHyzlsDqMYYCNTQjR/hrPvPykl75Iv
WEmTz05RsQ9qJT5G9ZyasgxzfEIQ11vX5HtOaqg8T+Sijsn856oNMZmm7TvKomAW+UK35rbpfNVo
zOdkMRhcQydWdBSciMfg/cotjcV2o2WJzMc6dPrGWH1BxBk9dhOLHzhCpktHUlc+5tn6FSbFk3u8
HV9E7K4W0SA4de5C2wCqRiAPqnZOMzQTUWvvLBmjT80yrbe5ADCvp5xHapvPqdo9Lgi3pMcIe3VW
d1+ostoRN20ckUCUKpZp5MT0lV6gECmjBdQlT051arma75n8/1q3xCxPLF3JkrCblisvxhMDTOGH
n4x/jsZc2NnLCV49Jr41OhnEJ7sImNxfn+B3X/q0lLWP+FUp3sIXtuib3V81J0e0KHwyF9jtnOqo
ORf6Z+2fqEeR40cWUknxSq2Ug5njzXMtNz4kBKRG/BmHImthcvTLvSZE0MiTilx8d5roWU8eipk0
1FHsD6xAmAPMTKr1JHgXe5bZ9tvgiWixskrnSJ2S31mhPzK7tDx+klrh0jf/2i9CHOHDSxLr8SeL
vwIORHXduuOLvkfzaB5VbRvKyewwh1u+/91cv12T4zq7r/EKew079WB82upuS0ctlzjU8qIZlbIX
K8+qa3dfP9mYv2qYjkgMxF7KkLjyu4ypQpwmQzMMGuTTMgVUJST4KUoy7IYJgCej9z8PnJC5bzrU
zUGQSPhCL8qCILm380Fqe++GlE1wDpKgWOJGnlbF7pQgrKc6syoLt8qPo/nSkgRzRsX8YwF/+PJB
aa/Dx4Zse8CQiQRg3lOJ+OacMc+sE7T9vnUf/ZePkmB0HcT8N1cIcIb6k/Tk/SE2ixVjNB2/Ug9y
SUqhWadBCDNPnIxniwPDlFEKaklrQryiOl6vyzdIGJwe8mbUlhQBFXVNsm7VrDpvTMEEW3U5yzd4
q0hcvRezPxGdL7DvmO2tXQOwyTafVi4A0sxLCHHxZN5GHt8cwNBvHjJZEmKVqJL8zlb7j1Z40Uex
5+EpoRVhFzmpEmdEvlEJMUH07rGTkalAvElwnvhmASyX8gy6UZa+UrtnBJ39fvTK7oE2YzJGy/o4
k7naS5VlJ+X12zZY6K5MVMa6+f8cisug7V34QzS8z5iroNNpjPS47xF3jdtA1e2EsnFDUPDgJVpu
dTd2uduFhq8d7HFgt4DFo/pWggP8rOJPGviVN20EbK4e6sTJZAy6yaAcL+hPsX0jz3+HK/NgQ5ad
Tz+r3ajjBGl+QLQLsbwd7xLRIWK/qGRPpjCZlTEyRGS7ZWj5aqyVcDNN3PjIz+flEdtae6vtaw6D
G7tDmJinn4QLOp2ugIUZBBLpqG621LM/DfpuU/Rl07n3VTS2spFOSKpv0BtbtckEr3obyr7CvZ7+
luiLh7W8JQyvatP3njDe5Z5p1DxJBy2rdJWCYxxOi28G2SePH3m/7P2QULMXqkHTz/moa1tTd28G
DFKztBE/G8309Xi0Snlfhv+LOvcmZEvtjbW6upIx6rh6ZNpDQCymDfciBGo4QbIik3/XnKdotX4q
Ea4ibwNXzKqDbYNnDfQOc0HHAhzeI9j1wyXyxw/pqNvzetB1dSbDX5736kRWDdTnknItJHKUzf9Z
gwwWjrgwi/ijaql90z8SUD2neFvw5qFpkGOYXf4xkwviseDLtKUN/aao4lIfLV3f/ucxuDhTrENZ
xsCf6fkRDV+qt9p/Tu8EoD+LpbAyHMHN306EEofBCYxBvodc9YqASQFIC5t4S5wM17y/z+FDKH+V
RnidMEIMjGY1ElOvWLVUrdd9GuG8r7qIboo4OnhZDDWMdJb+w9wP6zzlKYexpIvbyyqnbm4sQHSG
9TIXapVcQXoRxL640LqY20d1vuAJ+Htp4JbXXFdx/d5sPT2iUMFgboRMkugR4G0pc/Hz4Z7EeWNq
nhWALZy/iMygNbXg2K/hQYxvFeAxbDpRVyTD+kZC6XeoIwpZH5fOlVjhHGxIHricgaySi88S6w+W
e3MlqM6ya/8D1PuXDv12sAWL54FYlM7T3GL1gQAOcE2U+llbpHLw/5h87jeDUYevLQHkDlmHwgn1
JYYZGn+9Zu8nm3nkeCjEWbc8E+i7MDaN+ultIq7BKJgfwF2wdFl0YDdVDbf8TjXY5s7Qw3TGRqSO
B8HwodeAfCBYAHrcr3J1bk2eRL+Ix+bmALvIQDYqxgAK5ZW5U+Ed5DKwnUtpRuxkF67AzR1VxkHt
5rVtJwYmAbHBxHtrW805ZLnlfPvs7YQvx9ygBydK213JDfAnxWBycZtBbLS961K4ph9s7xTPkiDx
8ZLSDUA6NSNvhmij1BI9Gm1tw+XUCQ5lO7DqiY7wjagm5R3RRKk71+QezO7u7vhCQyEStt81rrHn
g3uYVXSZzSm0bi8x7eayZS/rAWrhlAtvEi0hOe+1N4gj9w/ODcBe2lSId88HBX8g6/CwgMPVJx0n
VQNNrNKtcc+xvzn6iJOZ8YCbr0pIKvBe0NuFZQNg7vr1a9VtboJarcUBIlHjVWhfVI9+rqNIhTtY
nM5UMyRexwM9SoCOkLzKGSX2JExCRtcWs5vfIuc5lS23nGsemlVPnwGmSCMlyBYlkJPQtfQswCXY
gQsjHFRzD1jquDt1pevdjfEnBem3hCbhj5dmnYlFSuaaYAeU1SR4adlqUYURTK27eZHkdAC/HVL7
C4s0RF4YMZshUWp+9vNtMa9OvidkPucIj0Zbs+aXNMgdUef4wYWyZvqz4kJ4Tjm2LOMfTsxaztEc
GZpJY/gPzfNlPMZ87pkaFEBNvLXYgNYIAoFmpkEDZsP/gA9LC+AotH7D0vrkxMXg5I7POSXCwHhq
YHXok0tgKg5MU0N4j8vmsvR3A5iPjJV9+Lg4Z2hhpylYcli3ds0CcvUhHUlt0cg+SKAP7u4Cv2gX
YE+vMjWZQwLPL9iby3f5ka83zexZPsenrU2Re8AH9gwOOi2A+C2864viS1T0bP/B2/dD3ajgGlCm
TY4EnFuvrhHUbK854MV9FK6tlFF7PuprWb0w30KyEkRY6ylcnRIUmfxW/UGaqDgjqqPpsvPNDhV8
7KQEJzgnnF22X+VuRHQR8wJotQbEAcF7Gk1U1N3fwfPsydssytNJ8KRk2K2iE4s/00HD7PTrBjDG
MxRuheDLpJZ07JAHAis9aNQxs/G38HSoRBTkQJCgPy5zR2dMNfDavsuLP9tmDQqdRoVvGrVVf1WW
ODxSo/cgK1+6GFTcdpDfLim6pRrliqxZgfvV5vorxPFk6EZFs9rpErK4GwaZlg601dNvSYlnF6en
2xQOQUCgI3vkiG662EGtlSAFzCqN+cIMnRDmX+QTNBYntepGpN9ysagLCi9T5pVw1GdWPExArOjP
V8z2I9ZfKlhNDbur77Brf70lbWzdU/F2mCd7sWiQGf9BguowOk0AzjwN/AY0uyc1B9y9oMi4e1kK
8AsoKWMQ6ZwqOMRfX9OVGpWGhRYhQK809O6NMT34alaRmLBNqLBwNEcJ+YxBA1j2NA1Yt1ZaLj/X
1+WjguhR5XHFuBOWj6E3mBL2W9yFICj6WlJ8FSR6v3vfxa7uWyCrdtujilUNXs1G4O2mouIC/1tr
MZ8DKZtRs+V8qHx4Y/9FD7wqt/b84rhMJKqGM77TUiBMwQTIM9HI3OFT0g7pBdpAFbUx479VGiBi
YiUnnMHHhtGyIFNzOXD9KYGev39TM6OslNySqwXrrdHvh8kcxzqxQRJxbPIOUND/RBXk6UaYWvKU
cPT4p35yTSawwhqW5VjvbsH3UAjtR6wQv5HSz2RI3ITeKZibv8H7fo+V0h4GmMoxBVeMlSeQ6Ho9
x6LEsj3kSDy8uJfUFNwHKABUYk/VzGWopWpVvp9w1iC006GDvHjEjIkBr7p5hBLNwpLDzt2xF27C
eOVAX68dqfKS0Cn0O6a/o7EkwmxYztBI2XZvdlAeo8Op6cT/mDu0KuwlT7pmItFzGS8DSFsWnPly
7+JdjegqtxyNnOf1VvN94r64iiyRxV0TdL1y+iwhXBrpX+NcJk04F8IheT8vhHDcwTwfN/WReRE7
OcPv40rJo8hlwPKV996Pd/xOlWf7RmzsBFi6Gc0T9R4w3iv6wggKpydGy5WosyewTsHaRLuPDr7D
U0W/fDXeiosru31cJ4aKXZYXWYjeHWE7GCDs9NckK4xlCfipdNbECMwBhm3S3td6cc54AIuovIe6
GQo0D6wBsHfd3xd6NdhXGRavtyV0dSpov7u8/IG4kDO0ICCsMAt8S4gZxQIpV8za8CudvfsDMrj/
lp9/c6uoWycKh9VsMxeYIFahz6yRviRPglXu29Hta0809Pzyyk7Y8rPTS6sv/vpW+jUD3tQo7q40
oXXKHEUSIpIKiu/4IiVB068/Lanv1vWBQWj6nvI4UZhIbqK9Ue1D/zLGDFECpPqorNAH1wnENZiF
2iIUfBb7iOEuVLMOOk/FTsTt/+ZXsrTJ2NlDD/G23bYFvnaM+1va9Q0IzhvvCg169917wCQD4cS1
0eOHaDNrgbjcbRmQRLWDLbYLwdy47fDdOPNq1nBkQ26OVojQBE8Kd3iND0T/w8gtuWCFnEn7pjM9
M4T/C7UFFjcZsZQ2wMkhOdVVU16gsFC9WDyrUB8s4TtktAK5LA/ttKfcyXnLZI1AfmfM0++qJX03
o+i9EjEkvj4OvFQ24nDMtZk3EvZ2pgW1hJdO+lVGAq2zwL9UgLpuEGGVb0jOAs2A+vodd1DQhVJ3
dZh2uWWx7cSiv7LgWk8rYr1Wn799KlzMcMiVs7Ju4z7XW2Uz/2dzldN89bFjiwoZ7kTS4b3t9AFv
U1HDGnotIe94ean49sBOYV1orukof+nf/ZVdBA21i8ACIB1XmWhqaqzYhRRGhCsD4l0e2m6kwM/W
Aiyp8bmzSdw065EmwpcDRXwnml3vSqgpYdf2qtls7EJBOg/vtSg9fw4eYZD4nDG1UNeTpj9xV1Nz
R/UqKh9bS/4oZT4jhjVVYNfLEuslyPXD5XoApGDnlH4oNHXXuhRgkcdgNf7amMSVU+JYFak3f65W
KmWkd7g8HAXkB1ZV16x3I4WJVd2F7z684weNKYRHJJDY+E2KqUPEYOnJLUS/cOB9iTPkt+RNT5Nn
yD+cKpRdi3BvNR2uZETyF1bMzITj2pWEmcRUyuvSdSkD2+69jkD67v/vHHFzLfNqEfwEhSMI19Pd
rvEoOJohXdOAWUCc2Bh5PY8W+uqVek7Cdox5fNv/0nptB7SbmKdWjEoXG3vVPtyfv+6JkueyiZRc
N2GD89FWhH1eBwF0J18vwO5RiaQ893OwkcJY2zBhmdD5xlbLycSPRmL9OHFsIICKA13fTxND3BRj
q9nnF0KSVbTlKj8V9jiN5slEb9/Mq4oIzKmVeJQ59PIK/DZMuBG9EI+hucKNE7tZbEh5Epl5wogE
q4oxOhuUCTjMC2LcO89SQq/PG9MULgp4pF5/CSB9wgLFvQlFbZ9ZuK90pTYOMMaqxXYRDbSH74s7
pImKf61SvbR44+sAkZ3YFEpjABOpPARLzazDRgFi6ALG7UEt7TlhafJF8HfmRL4fu6mmtUl2OIWS
8iIE8Q/8pYMflNvHGqkf4vOZZkYHOfdeckFItzGasXf6WqwvnipgxehafJaDxKGq1vwOnmtBZZu8
s5eHjXzTPV7vJiFey1obP74JuSmBV3O0KYjHdCjj0O14A8BLVPXaXETOdktHfYC/iSqHjDdm0hkk
GeP43Sq5ysWTaBUDrnXJk8UO43mfTNi15vt7tw+JDazBUUazt5h+k7mVC+II5BFnEUNHLou89m5j
yNaYWuO8oXUhT7CVSc0p9I1P8Dc+ls78NX/4jRZtrr4IySa4sic6a80Z42nHAGDGqtHMzF4RwSLM
dM5RHR4LCPTN1Ps1m9sNLJUtxIAaM8Qk1MOGGCJwTIZccytsRSs08WdSrTDO6bVRNp1ieoFd3Ywz
C78ThpqzVbehQvLmDDJQPmy8rUjlFFeqsDALTkdxpyXc9ZZ0nVKleN53iok56JqEujgWKlWtTui2
LUPE00qMipEggXs4UWSFNY0gOPyDNA7/q+AUGT1uMJWzzr3jKM/T0jXMz8MJUQTNg9TNsw/Cklv5
jg8T55eAGXfVkZIyuX5Y9pkrTZr4PTgKt6seOa2pKnVHiGIhLa6Qs1NkSJpaz5J5crHGW82o4ekA
bTaIroutgNhbUrcwnmKLsr1jQAjY0bzM9aEenPvTwaSeNGvZzlsw4ycKPlhD7+YFA/sfuPDDVSPU
ILFfeeSiPguxPDk7yYEP2AvuD4ysvopEgv85QNxPz0vkOgSv5bR9pH5WUlIzCHu72ykkS2Hs8V+X
gFAKS4dOTrK/bdZ2Ia/I8kmh16IxrDDHCcv2QUScqXHlOEcDNMK+shXULCQYNk+YDdK0Mvs3CJZ3
XyugiaGWRxcnmGraTZk9AjurpIOmXRypwW/lp97P/FdDpg/vYjXJw4XeEmCZPuoabENnKTD4prxs
55Lw20MrPBwDNgrWo8pUvhTCnhlO+2IX812/bNC9qCHtCnNpH3ydEvsmwVqpH/nhZUXFGh4cvJaZ
QT4XNMI+dYCwKysR1RVqZwUkt8u88wDo7ZbNcGgQLS2f7Zr92nqVsv/g3Pp6ywX7vHFkZRzqLSeB
4E9+EzxYL+mtuHAoVRcjWs6QXjLxN2RPn57nfa9dDlcUjF9hvNxPBCyIUr6IcHTMJ99ax2TV4NTV
poAuteVZQqOt6k89bhjyw+DB0qBDIfhnOaTp5kUXpJglCBOgWbthHYIQcKw3aXGeu5KowVjOXE2B
nOuCzhAkG+tCHSSiDE4SkK4NlcLXbFeowh6tn2PkKE+VuAhw7DNXryldqPxmqiEZamg0uMq0Zwqi
fAJKpKji9oIQbKWeZYD0CiLw5F9ndAPLU+VMAwMTavAQkqGA6b9sf15LFIsF1M6zEtaKsVzop+O4
PDIPzgbW3kuxZb+mro0veS0wB7Q/D5xK+LVXFPR0W+odQfxddMP1JpaCAdLl/gIJ+L699QeOB2GD
ttOcQvlzUVk6S8lRoYXsd934GSyCgYgTWJwl2PCu7V2ll6skR3gro+JMZU0cK3Sc3tqPn5QWW9GF
MEmIIAGdcpYT1lLo4H1+45CIhd8stSjRDqdu4SzTprGlT2GJu0Q3pr/eKeg1MzRR0yilyGhQFw7D
yzv1LpfAY3D3sF9wMbQIep2ACLOWTjuG+S3k7Zvhkbpv4YNqXY26zInB77LeDuKrTGBzEzSFsLfe
DsyWHGYSkaScUtvlaUmCvP/1owqtJdur+BZzfh5yg3wyy12UnN0j9dz3ce4ESJC8yYdQD7nPlHwz
VdnIaUBSOQ2zl361W65kI8CAqZ6whO/7Dbwp0UzdmHg07w2R8bLFPgRO9bEgMiqfFGX2OiQ4O/gp
g/ZokAnKIcD35nhjWbDkr1v1/Q9rEPmWOH18amJDLEpXDtWX3eAYbSwr+S8RJISn3HlV/zOHNMGw
qBSl4uTLbHJnv3yFWsQAvHuIqKwwb9m+Hkw/t2rudVFfA0y/cqv4NrZx17O7KEm4dHraMFOUdPBQ
dnluu1k8rDzbO3ra0iWVzrbDpEilI87+WCo2KnZ2Mfjj1o0kWVxylpDCB6EOFu3cIa4YrKqBnEcA
Wm4gaxYeTl7W4bhx+mNCqF4jzpHNQvoIqex4H1TryEvU7LYPkl1thSc0zrZaurYrnXBZzY4JF1SU
HtAb7GyS6YuO6kxqLO+D4Jy4egi3QeW8nqV9OlsU/+uJ+NApuQ1wPIvfyk6KUfq0IHWNQsCmziMS
mwYMtcgDibe4T+q/FmtIw0CmaIQIAuFoQ23rpaMkSxGxNwRS+hudGxqBtec6a7Us7aKISoRShwM3
GivfaOy2puHuQxNrfJzIKwO6Iftjzf1LAXN5+Nrc5pBzQmK2eVwfA3EoUXr+eu+ghUR0NUdb+ygm
kE3d7Cm7rDzHxV2AQAJO7wtg2b+WymcfLBPpTUvLgwuvV/6a3JSsXT8zCcnFTkINj95X4D9a5MJK
knctLXd0dl9fWqUmms+nbYGGMUVdlPAENNfzarS5SsYNYl6rc5oTq4r4k9iisq1Gd+vN/srjlTC3
U7yYncIwxF7Kkw6QpHg3SYdrY0NZl+nP71lyCK1JHP8V13F8KrXK0nW4tlVqeLREJpMgjMsJxVUB
HelthCbDsnyPopMXnmVCeyfGpJsCSqq0C/P8tI5cbGcCrtAA+yfYt5rK0ErQdF8MWwwN7t/YbOEX
crMRm9/vmKgfHRWWdsAdo7dS9x8p7OLQ9Qno/6ujQpf/d8khQAlA9m9kO77G6hAh4skGSaXXdhjV
6ZQuQcqmt/7dmX28q1nPKuN4Jgt2H/AahsG2fH4bVBbiswW4R2Ys3Wy3ITyvRzGK+ZZYzUqSJDvV
p2lpt8fomg7cPKYbytzV9090yVmjNRvH3qbhV5ErIDAwQs1Rk241Ru2pbE7cSJD+WM3fSg+4c5Zb
Cu72z2bPM4hBJVJEit1UC+hPRHquDL1/UD0oEIujpTe/We3L6Z3R6UPnNP+Lty7HHqr400k1CZyw
95cQvN+6TZwKGqC+V9M0GT7tiYQsR+AXvWuh0kza40f8AR2EDQkOUeNXb76cxOS3BmXquir+gse/
lK7dg4FYKIoIGg/aMuG2tHmTful3k04GpILK3j2yJOnfvELSGwJntepxSgLREznzQXqGDUWc/yxA
c3D8yCBbK/kRvsHPdtaBNCGvikZvBoMbt8t32mP9n6DyAHcM8qUD3DSfHouWGgl8SGi4dfF9lUmM
hzhnk63HOq90stw1PzbzElyvVgOVLYtMufzh8pdm3qYxvvEz6wTG+p1EAZV+5bxGsIIbaQ/kqZdv
G2MrmKxm+JnwSG4Emu9ukzZG6vwLTPWS1T//kw+rAbs6uDuWry/0Cz14Lqd+0RKYV1/+3FpJh90u
AX6++7ej29GoOf7fp3k1hzVQF4cKUuBqV7uiQvUEHk3QmLEEU5R6Yh/dFLmYt5YjZEtleRBM1xf1
5j03sAxJPM0K5omUMRciatL7MeqUO2mr9QxJnWeTw+fmyNJdVNuRTzUkdp4DFaSaJnxo2xmSPpEG
Gp/UiuSHHXNh/u2xGjbkJxTSy/VkkrfQkdbZgrAG3J50ZKF4k6NktjLVOwqJXAwFCk97Ub3jIAWs
OdptVa73dT6720A7UfNI80LFwaz3ok2En2KVIc21qi6KljIGiw+GjydXbTWNchabTTITBuSPwVMY
lApDAhQCFqouQ3HCWP0m/G3g5Wp61DAvKcDOf4wfpIp+72eSyOoWvjV5/q9LxLXPk5bA03G4gPE8
BY16HZ9OmZKMaqHMx0q1V3YsRcDiX1/QIgc4b2vQg9aqmOT/lE5oEawXfCbrOZ8xhAZACrxLT4Ds
jpQs1q7MbmHXQi/NXVYZEbmY6/uG0Lcc7572WKAjuDbwP7PFWfSCvjwQNRY3gvr8OVdHWFw86aTb
k+9Sh0BKS+4TlYtyI4p1oKojm6125Bo+RajQsnITD8sKgdlFvTFqTj1nStSSwsckzqgsBtas1HGW
w5+I7onLPU3vZ5sgZRdx2OpSTMz3snX83MWagLzgpWQa7t1fSDsOIkp8XgVWkRwUpxKua0A7xd20
L/Zjd11xsOiOKYyK6F/V63SR+VogAkYK5akJop0fnFdV5gpc+ioo99Tsf+q74eoeBBh/q4/r9xoa
wI5tQ3QyN4UKLsr2kU0QvxrYLfjLolpNr4ZFnF8eTybXPMKq7n/vn6vuSuImMepy/AhkEDRAfEV6
inOkmp9H+IZP+8PTcd3YsBonpiEIUgFF5wVc4wDVZ6PBveFvHXuF+mF35NSXh5jhs0KTL1Tzy1b4
DFJNvUljaeQDFpMl/2CjiiS4FI6/B/V6oRF5XfzSmDEtttSzonL9ZDRFn+V9hjKLTg3C0jGJ06C0
ZW6ItgGcz3o9LkHR5cboWLKOx3OG2s77PkiT/N3jt7A1mf9cyjdUoF7DmFoAf8Lg7EwdefdXF+co
0otz/iyYMLlqZnNi21pOfibxAbfuPx1p+KT0CUwwgwXItOtKg5v98DqtxIr738jsYHs0P5tEGfyl
U7XV5HcYVhMbdwoSvyLQEE8icOaQxUTi+T461bekglibGblMTAf9Gji8tAK2B1exFHmfhGooLgAl
Zhz+Uk24keYXV6v51H2tkRJYdj5xuknACRWdHEVlY/7dH4LljSY+zxpMJ8s1rqH92qeplxis/Gow
NgTCSFRdBA8hu8UA24KSvItfN9qzOvVRlRwO8wWL6C1v29kTyYg7ziMuWANu74wDaeqGIcMWqyBS
0A73Ng//m7j1ZRLccmmHzyYzZpJttuJ36yA8kKFBauQ2l0Kdkw6xy28gJML+7hzRUHueK52flbvh
a3dAkk77GPXzOFXnxyaG9R7DcUH0DNOtb7SjwkwX7pdW+Fsrpgz+/fZeMeWKN8hlx4FK+MroTvHV
lA3gj0uCha5mASOO1LLTlIFHT8b0058ILK0wDRr55z582kWchNeeIcftKbS4yiZzERFqLqM/1P5Y
2gvTFpSPd9rzy7q6vJoFpUICRwvT23gw7lkvzOKBJ3T08mK+sU/xQ7kcRqhG+CH3PTyLlmJzPngf
QX0F3pAZowGMdz3qggGYirPVoNspB8ysupMf8JYV1GEuMqJ7Zb55jETD5oFe5keL+h8JhaWJJadd
q+pLkY/ppumJGJe/dFP/EKSg3OZnEtNVtQMyGohll6sd1Cjn6bESHtNSt1bjaHaYI9/6Txg/h8iJ
0dDK6RxeHMCBnzdBG195iPi6n9ZHjEWiMPFYHba2V3v3c6YL+Gm0fOGjOxrEP+CXc5YB3It1Pw6c
wdKfptQ0I01fWqVyNv57+APeN7SaT/kTDdoMIFBYB893GqBwikE+9UQvMkizeheoQDyXSIQXTubO
DbqP6tc7tmTkkxJO3aBc4U5Em6MuEXwUOrxt6xKCrsEatvEJaPG8UBKxeTioJEn2/A7/K481O5XV
STgLxGEMWNctfV9BNd3XKDQuyCg99wro/JwrCyMCSKh8OoNzJu0RDYOQFPI1iF4M5ChBJ21qVriw
ZJ4SynWeeDl6thXPEQlZttBhraPfIOU5MCStEz63g7xbo4JTAiZcIpRCChMxwyn/2mfFFoGHwgmz
p/f3hzrcdKkSMyxyWBDabqnaYXENNDVIbbhcH2/5aLB8neEWPLnUiGhjchL132yZeqAsDsXhMOzj
ESd65piAQhp0ajxdttFDsBQ2inHK9Syr16S6+fRFQC/fTE3/CwiVc45/53eOZZhKFyTX4pcmhmgj
1JeLeZFJUSjFPGJeiJVxReSqHBSyVdHGp4B1K+hN308/hUc/xgwrGVIf9DOfpM5476GDyoHfzasy
7UmP0yrXb1jfJsfq3nxWk1OcaMs40qC/ynXefFcDgmWMUb7DJ/auSP0wlRmrXCbpv3Wnjv4TOMyM
ogtyY0AGJPsziXOdz9Cj/9lsaoa888P7mEyO2ix2qSPm3kymZMQxoiSPrSgMiaz/r4z7bYOCjLV4
S9tGJ86iJljZyCp2Ne2rKQ2qv7fXZTAWj22e3Y9XVW5SMuirdln613qHeeKlNBncjl6g5zuzOc7F
5FpUZnRKqURbQxzXCbICfbmaFa3wNUmpQbrz6YCIKpE7wvTCGIg5Nt4lXyeaxsGOcaokTNCg99wF
2Usc9Jnf3knos+nr+ndfM4gZ1WPm20uGY6ftt/RlVjpbRLiIZqsbPZokRvhHzyWnUrJOgxpEEKn+
JnEKKlWeZkIm78YDKchSH5eJORj725gNILuAKDWfXoeOdYhgPNhU3wj2jyK0y3TkzrZGSmvsDmfY
oD5SO1RmHd2HDF2hCK03ToMKlsXNekseC0unDt+VXFzQMujzHJBQ0v8mXmBHpXBMx6I6RuQ3q9s/
2cw73j0m1OVCrOgCjz/lk0M2cpcwVpF4RQ3D3rSpMkCJbpb1ijeqbHquy5UZaH2AxINDCkt+h0e7
6SsiilPmoSmr2yc/d2CzrXRPeRYMbCqk1hCB/eoPVABiSZ++gepHHDjFyLUEnEJH7gX7Ze/Sq4M4
WYHCyb/GNBPvmfqqxKGH6dCpPsrbgHeHOz669HM4IWeMvCB2iix9Pk0nkJnsz5+NeJlnVzXx0Nvk
3LEdtpSda4SDjY6AQbmLEgxwpqi4UUhwfqCcq1ipGKOXNo5aeQ/U+NSfyvnVaqZ4grmckoZ8+WVd
UTayLdc8XqwqWqsaXubqWhkpm6XGd1T/KMAjGP2z3p/swAoq31y0Sk0qnl408Vv4bCY0P4HRvsSR
y3q/EHAcNGZFaSDOpcD7LJ5CQlDy5O+3J6OcPqxHm9hnw/3ATYHXs08x05cmCQgF+rLCu8E4AVjt
SS6sE8Xz4McI8I1j3msxpBUvRv/tMkPJumRet2R6IbfHm5vuKI79cgD4QC5e4Y/vqJxuBUZ8TQxJ
6nj+lbxXno7EGHLS904AVWMrzGVFSxxKK92frg7nMS7z3Ly2VOnDo/w3J+Uto7MdD5qboobExYF5
Y5pmZKUEWbGZj5RhhWlrnAN21hVwDNMw6Y/LS8hHPhohJ2BvBEeVHUfikvwajfhdbJks0m4KWuvt
J6tmpsxNXECOeTdV5+lN0XM9crB8qVN/cLPTBqZYxsMklrBDAEd90Ki7frz6vmTeXajXRc9ELxpd
IvYxBBMwh4sK8TEKGrFnXgpb0XB2XjBskLTMEWVSO9mFvqBA/rNszHU8sLrBPAMa9X7ouHBS5Fsx
gP8Zd/1IyNc4PRmjk7aMMyEPzgMupfjM4fec4lK4aaD7LrvmIsPweyaBjenxVMqYuXjjvaa7kiVC
WvLAr1PERdvbafCck0IqU9CaFW9/+wvk7vAD/uKCRjhu83DsNGE9Bbqo9WSjzCW2wmnDpmg+EFGV
Ot3KuMvHb6PsfzQoxVa2RzhOQ80UtToN8OPzd1WK8k7uhRkFw2tgNeRFAjGsUyVgq/ql4m65XOGw
V4w91oozcq2bNdfC7dFmJBCKUGL8pPaSNcKVVow4Hk598GBUBnBlrmKFE9yxMHvwuqh8X6AV8mYU
Ens0oLXrkklrqgL/TJyk32eV2CKdkdVUBXvpD+HjmXnudVhoZP8MIcWmpSL9L7cRliCsUp8rovR8
5D5vloU8vHeNLz5jnl7lqE+H5RqJJPFPspyvJTcRWEysWOEefdM9V4616s1N6NX3jLr+nZ+6duOn
7Jpyl9LmszcxFhUl1RHtyZqSqiJtn8XCK9nBPvwb1GzBAeaAvmxPDU5pfj33psI6s+X/XaW8jkBg
71JGfvrDdgt1s/bf2JqEoxtLVsQk55J5hAvKvENFizmlxBoapP4HB7/rVJC3uj3py6Jy69VJKLP0
rR3dNHPIShlPKQ8RsxGPgSvVFh4//TyaJ2SBrLgffcVPhC0nOSE2YTXaiMdqfo4LY71QROM7bSm9
cYCN9s8CherEnacioDMKlPSCZaLQtnojxZF1GbMSQ09Kuv56z9SmFWqw5Qebl+zwQWdCjEO93eSL
I8qndg3rBwh30GiM9VzGGoh5BKqnPPixoz7XisK75LiS9VhuueTEGOjdWFsfEbkwHpRRIcUp6yrh
mz2UQNAjdY9Yk3Un7VHkEY1emzAapHZq4ZG9I8NyZtgmAxDd4cGEXmFPmzzLPqBiMz+8pWMq2srw
qk/OLMwxmS/Tj+NIOVlSmSPKBKiIenqRRdQNBQHnKeXDyMcddi9DdAOmrgw/V6TLViM4stZh6CEF
Q5oVn2mxsO5V1OKhm7WxE6pHM1sg6Kbz8SxYfaBhfOWscgcO5FQJ1Nusosap1pW+AxfU3oz76MR9
5EExkNQD51T/3RM2EyWlFbq/kLVAc2T7gBbyx85XExYj5kjpqe2kBGtsS5HxerfPD3uYXmFjDNGc
kUZp30Z+Xz8MzzKFxg1gBEt7vBDdkB7fTPezV9olSDeo/PqfAMFbCnvdhdKQpxzJRDbsp6wVSlcd
dLyfAjaL03Mj8CLVye7xR4Q/u2IZ9bpYATHUG4MoRE8f258ckiTK9aB9RswWv3B0dRPUiXPzREd/
mgOvDz/NZezRjihVVk/ivM21R+WTCo+MymlctaGJj74P7BkkBsClA2abWE1bX1Qdtqsule4N1z1u
styllKR6DMzxvfuBXsUM4HRqMQvsAJLK6OCmHjqm2ZIJ9h+K7gunimOc2cDge9oN86vwiCfda3jf
8qZkLnnutKeZzoK0Hkz6aHMcS0NewS4RfRcUSXJvm6xiA8aXcnj80iyUYPXsK3rsCitNBt+30M2y
aICqdIhy6kM4Y6QfhOQ00OyyXx9mfkb7LYd5rUXssycD5umcylFeBFAklZyNITw3J1/F5cQa2jCL
lwR0h22+mnlozKKo9z0oJkuwW88OnyiJN7GxA3h2x0QoX3daziwfUpbTZAjBNdlmAt/4+UIP07Eh
GkV4P7OACmHxZgrD3yBPl4HtNCkDbN7uAK8LmURKNjNPD9Xlowr+B3PtSdF2+MEcbEyygz6VWrBV
dYmMM+TTJkPPYC41h305SAH+CHPbbNoWej9Ds7m+m13mgqWQRHghyikMI6G+Vp3Psnd4c4P8ykjc
QiIinYDcuH6WNNYpvWz5dkT1yBsSW1Gk+fsLkPnckGblx2KlSDQUrAJjnXHPUB/VQUXQg1Gw/qMg
2PwkQkWnG9+q1MGmlVY9yG2tPQ8z4+7XHME5RmGvzEgjQGeuEPcDUX6+wCIe6tS0aSG6HeKCZs02
v50nzfslWnMQE4t0xDlsDfC+0pHv/PPYGt1Ciqur5pmnDGf/IC/TSuxMay9kOVeudOxOnPewk3j+
IwMMdCNNHt3osLQ6pnwKvm37cWSpuFqyVXRVtioyHHmR+gPLQPIJZWHgJpS2rrSZ31JhxFeTjc8a
NANZpVJNGMNktvRAhip8ZJDU+BtKhqIypcjY5p/gPJ/W5pE20MlHr1bA3ziFS0zWoa5r634esS9k
V141VD3iUa32RaSdlQAAlEhUrdWmusG/HYTWKTaP6HtHRF+I7CAfx/qiMqhbG/tVqAxRVkIa7n6E
NqCJRBg4Mq7TIryZINQVyxh4wzQ0XBWATCLR1N8/XyZu3tguOw5dq9YFS+Klu0KdnbrYA4pDvqao
FghAnVqfykURRERILJXFvifF1yMqHjLr1jna9Ay+EIaJ3hAY/D88BGFxzelxosbNyOw5+U92e2wd
7FbUY59WzGVfXtJE0qMCmyMVp3z4XH/3G1UVGA8dmQSEflUL5jPZ8yIV+ynsU7rOT/qiz+fn+UHp
shNSp/U4q5ZkO4S7vV9gkqvIEfHIdnKhadmO8z6XeIhCOg==
`pragma protect end_protected
