// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HpE7GmGQp8XiVN8V9qu+vnnRcFBuRDUqxPeKTebBs6zdf6xVZ/UU/WW7aQTd6UZ1
8IOx1Az5oPsNNtOZA5dSsA1xggWM77Ef/3XrGvUDN6qnDhyKpKc82FcyTMdnQAc0
Pvh4OWXHi2GnGwFSFukMfFrVX0fFIO3uzjry8ovJFVxJ8jf+2ojNqA==
//pragma protect end_key_block
//pragma protect digest_block
LlDpTSDxKGquahXaqxP6oBMSzTw=
//pragma protect end_digest_block
//pragma protect data_block
rLo9jJD9Kf4PdbeWrcne3ecae+tPuSs3DtLtdF/GJp5uXqEpe9nap0KkuoOgVz0F
HKz7c3WDwxBqRU3C0GNEwcuKqvNSA4AmdbHAp5m8211kgJw5bIgJuW7f36bxsObj
8CeemhLW9u8nY6WpKO/UYLipBGrnP44I9MMD9EDelfG8bnRi5L+5C6MuNPNAkld+
lVIEtCYaSYzfv1QaWVn+yyBEfSJI2sUMF8uJLI1TbuuxRzL3cxJbRppYBZHhgxND
YIROxfsZF8ST0ht5SXLTfgqimOckKqvjB97pSBsvkq5+bdWOvkC2gDe/ljiXoXkI
ATNBNZS/A2qgodb2uyLWoz8Gri+Pew0cr7s/3wSEzjnxPi7JKRzyA+4P8ru3cPVe
4X8cJjfh5MOWgn9MOXfy2UJNvtGTT0Xbvv/DPxbmxQbGJN4fwKKZgDWAjqL22uxL
owvq4vllEW7vrvna7aqBtze0MItLnuEZFWDanpbmn8Em9C1oTaGzKYknC0UAVzF3
bk4yMn+cBj0Ndu3Y3AVLKQKI+p3B+zOhRmPIlMOPzpck27bEC9Qd4xzE3O8gKJtO
kKFpTzLMPn5kqHtl1O7NzKjcUU8gxIDu7R/nmAWsV0jk1ZQDQvLgN67+D+pvSyg3
STGvDYwlCX2pLTC5ELcd9fRMsC3isa/zr4I1fTbobyV1ffzQETjVWJDUbxd6y1ti
bI/V4MEc6JxqpGrZWVKD/OIZ6YuJ0f0nuDfgeO/O9qYhayGfAdY8Pt+9xiA+l/Td
lyOX+M6KSREjN8PRYwbzcMFTlEfyYdG2H1/JgtA9l1rylH/7o7TB4Ow0cPUo/BWV
Vi7MLY3YvIPbAGRjpbd8FMQHFHVlW5da1Vv+quvx9GnFPSkhbIqeG1kDY0E7ZGxE
IsndG5umh9HnLgu1Gsrk2h74l3XkfwqRdJELeQLckfeZvN4xJ0y+Q7iqNQGKlO+w
AiYvw4DndDFHHXL2Z36GwAHK+MYpq4IaYIFHExxCKdJ+LtNJ1/mQKaIfgZgdtFpR
fIhe/HGnaVFrRiobfWiZeBFvwtHu2qogs9GOBmFrCYrXYWpMWKJe6jKL0zfUIPAR
N8xWU5kIfWbVXUqDk1o4WJHOFi4+JOzG7e5FjBYrwhu/GON+z47Erbe8JeIRABH0
BJuy2RwtU+Qc3v5ba0IMx7rDVCNuyg0BgIkvbzo6xEiGPqffx1GKSJ5aHeCfuerj
AeXBE9U4ZeKU4FAkgxq+6d0ByyY405ULFPyKZKmFqY2UFKbS43w0JxJMVpYxiOZd
IWJKBlE7aLIoR2AX68nlJZU9ZbohDnBP3ICENORcuC2DAhjOb17jrtpIO6cOYKpb
QicqPhRiVVd+GcluKzt/kkdlOQZPtx92p7r5GAGxg06P3V4eeNikrygUnl/3eYWn
fCQl3VqEKOi2PsU7ujDqQc5dd3/A5XtCKdJ98VKB61H+QxewEJ++1nxp/pm9JJUT
NQFKW5cVVV+kb6+Iur1MEQykRLwkG35sLaNzUtht6GapWFJVP4smuXHnxob1wT58
Kk1duawrXbolURo+iMNh1srjq+XBtTIZzc5uk321JHJnqY+jWdKoAtk8bGWJ9GrY
JqRY9N6O7Wjws2Xdeb/JnoqcbKHcX9ZQ7cTZq2zo+vgFQjPkpmX9KZyylD8/BqvB
5LVjqArhNFaFiiFxVrpTD1esndzWK+OO3Fzgr28IlD3s7hoUDIpdFC9cFju+UelZ
QFVWBK4kC38Zj0/KqFbcbSK3vWT/jJl4BRFTA9ijbknx5RpVBraW5vzG2BRH+laW
dHR7ciiDOOvx1KwUfINPSKDAPF4MsUtyMZ6RpOrKRLZNZbJJeZoTvOxrONMcdkWf
B2PHK5ZBTB8x4MUebgzp2JP572oADcAgpitetlPeDbv3wwHzGr/sDUVtmvgLk6vs
PwatlJ6MqBIDupq1nhGJQrsMGhXi4LG05CkOWJ6DoZunFHFfItTW0t7YosFBkGcG
a5Aq5MCS5yEc1ikCP8jg1Kj8tYvA6YT9rmGFdVPu0tniISZMuKqhrqYGWgzNVFP6
MuJYK4c6FUXxCOfrYw2SlAjkbAZoIHnWo0286G9cYLEtcokndN9qKBTI869fl1+W
yl7pe7aj9XDIqJlobW9qvF20ySy/L1HCfZ+q5cDd8rMRaIVCgjpJ3UVJw/Uy9Uix
ggYMdcmCNtcDmAlRS23OsejSriyVPeM9zLZ8QppBPfQ9L80AO4wiaCYWDDnzs5oE
bDCRSI7e6jmHMvPv/8G8o0IO4TbptsQv0Zc7eyAwCtaomGlilvP+rWUhDPZ8isEc
6qYm3Jlm0JJhPdfl4SuIZ1UnoPDPwYzZl/CloEZq0jRxqSceonUb1dS+0lhpIFy/
8q6nQJImRe2zQYPDJ2I46RKEy1B3ilaFSKSFLLmaxQirfDc/gtPK4q+/N3lYkvOX
NiK9Y82ti0R1n5XvHeavIZEPDiKDOd+r7zjv6H8DYUvMO4+QVjmnBDd8bUyx20Hs
lXb8qplszeaiMZo3QjXG/Blrh0xD5lGmTpsJ3yhjU7zLcNlFvBgmDtwUHeYq5E2o
rg2F6l2rfxXvGvpjBWI6e2sxI9S3mCSBPDTVJyZGXlji8X9du93Vkii6R7wIlbSk
RI1Jw5Lvx65/w1amCNlV18vJwQUB3y35pZSVKvJbq43XsoZiJ95y0dJeYCj31NiP
HTJMro/WJihqsPDebyADZC2rxaH1e1x8MmwosgDJKXUbMaLDnG84LEmY2yfQ5ahS
fvs6Gfr7m/cyHqWr5FjrrlqXhEOa5SwHi5Q4h1WYyXja7vhhe/EUcw3FVrYcRt9M
RdXSlH0tdewkJ1qAoShXnDTSesfmzS5iT/gAPemF7CWd2ooL690h/y2nN0HXFATb
TatM7BcefjUfQmxNS3FM5g+5n08pk3EtdK28/ssYavZUijYbiqM0Dz0hPklquwh2
I0Pu8aLpL1HE2mc1AefA+JXRg0wIJikFRk1shsrupXrUquczpTE8TJYbCX017d2j
qvUZoL9RP3BS2ObYt3oeX7Mn6bOQD8/8kOcHWP7zbpBbPbSpeoqwHpzPTBoEXuuk
yVpzHfIppo+IGUrbg/eodnTepMghW05rmZgyJT7mdJRgj3IGNgZ4ktsQoiEmFlDA
eY3fe+PaEZ6XEAPGIlx+JY0GjTiF7WoxaP9tsrVU7VdDwndspixdOMzTsYKORhJT
vqsEr8JtYJdJqmS2dtsD9BHv92eyVXc/tTqZgpVkVqMJljXT5ghHtJIBfIg6ulwn
P+bflZXPyGSrMNuAJfSNFsYYzMUBlAuApsZ6pmymLElsQL2+c0/I+YvD5xRxTbi/
R/5p+mYJZ7wJDnNnZDu5oPSv+JqfFMJPthuDF2JP6MaxdxJAKzFhpKBPP1ahswXR
WH4Qo3sHlPOTlac20PKi1/owwaRm/fdTvq/GRoOw0qQuS4quduIDoAgf6BTp9Ud1
+nKWIAMuHut3RBrmVS3ao4Kw1XAP+aWzUYRr051pBzh/LfBljcS3XtxJQ2Ge1iwD
rF8Q5bT/YEHAZJa6uqpSAbRvytJHFVVBW3KeHTbsOH0EHSQmNHhwdItkfjXTKKVM
GrzwxHoE3UK8NwfaGLFO8UdGPgOu+QFPAeox3u5730sAqgUUYyZAHTI5r3IuRQX4
vjyeatrygv/as2OXYVqZNTJdz3MzOIaiUDs96+1xDsm3KF/W4OhM81HGRQvv9wGe
dCLUY6rGqS+yfY6hBC7I4O8ZmBtQ33kbRHpSNAMhvx0OuG8A8u8N1mFq7GlpLb5x
Ko3WvSdYY16Q3K++RtqdGu6JISdav2RxYQKj/f43JF1HDUnAp+6u/dPvcKxlTqER
PUZVagzNMnanskO7anvHyFBm4yTSPXKb00z9a7MRWINHtILMtXs5MSO2eEV0THZD
hMeQqCHO17HGRFtIGzlTk8hH87HjKLEMObOZaYXPlEZUWZIRiA1gF4yLqTPbKo+9
AIPUxt8sblGJUlZB6u6OqD74Vt0+h8otNyjp73jXDgc1UupbTDTj6eqjdE1317ke
KWFunx7uSk7IHNoy3tYqWLyiD7MNS2PiHfpoXNFqXHO/YeuGev2EV5Jzeuzof6id
1vB3LRlbTf2W9nCkmL8sSpCMMTfRCA7E/b89qkOqs+G4GxMqKv3zWPJ1AiLechJl
6KLwH5mnQoUWT9dywZYaawQ3Na+QamnoGgUKhpRQdEfSnz8WMVAnS8tQTu70MVGV
bDcfdncNkAr5nywtKkD/yD1q6QKZUDEOyHwGN7gGiLRz2ok1elFjLwjvJFZc764z
wGeUufdeRl4kHcYbqPDn09AMtaRQfvGNHxx+MivLZJRW4OozrEeLexTXHil7aKiP
Vhi7Je/XSM7e9idWkTEmKmDLuYqgARccve0RKab16qSkTdhLgn0lV4fyHz6gAePe
mDSa4bslh2ly3tzRozK3DMQEbqf5syFEg2zDIN59+umGvLa5KOuHViXfEwuioDHF
xjNqYsdLCNjnjb8S9naBNMrbKk5ERLlL/ThkB97dtEj1006qU9/6ZFZiEAafUq1h
5q0AnOkZyXQflasR9vQ2qDE7/ZOImj7AsXRtYPgZJW/ImSCumYX5lwrwd/FrJFrP
PQL+l5HxcJffUQ7OzeDsjSha7xz3+nCUN0jeK52I3q/kN/olmDNnW6iaeySwzsb6
HCL1oXsGEOmIpvtjz165vcO0WFBY0xzhj778EDJvxYVkse/7dhC7JctPcpIwQ7jJ
T0weJ1jKHELD+9U610tuyhmlW39eVhjHHHvtyxMqL/fOZLPwnIceI03ABQrUPSAf
NTEd7KOxgFBdnhXsK6HPsbo4ZSgqU6hmHDvd23j9S8EFxIxoxDKbRErp4C8RonQN
McUCLU3ipSDkkHOTTXzfv008D4Lf+XqoUcqNfK8rT6U5cN5R5oIXdq9urTGRymmR
MGV4PYDs99BX1FEzS2reHrs15MWf3vzObclaMvsiRPHwQbbo5jT6um6jx1dmP95V
NjOQFIpMpK1E7RsEMTeURLmZiP7UceGCMYBSo7y39kiRsFGJhPc7qs9MAcst5ju8
//XlBgP1SO/vXfiooln4KAWfRzWlbdrrqazg42pCWAsndxVnZ2K+5iYmc+KDcdWm
aCEBS57yP9oTQ8tW4aCD3NcvBPBw0XyeEXKnvHaNJBkZbY10+MVXw/DhYNnwyYHk
qtTPvw3io8ivNl2dDkdUZpF3VcCMLPKJnyx5x2nUXMH8bRqiqSdZeXqairU9ydRh
VtyPwP53nAP0BQqQkQoDW4msuXv2upUo40OGXzHjVsdRkc7NhhtMJ9I+gMMLzC+R
PgR3iaBRligT2Z2PLO3ls+VjgdPvWM5WgdGzHPYXEaTr4z+m0omoFMN4iLpnuVoz
JByymabHAP4v5I0ViIj3Xq7CTke2bifia3+ho85fiwgqWxjirRMBxjp5st8YO81B
BdTCTm51lzrtgB1kBMysUGeFgfpau05G24EMOpw36J2VMvZLmJ2LVD5DfLvC+pl3
pDxaotOdX7l1LBoTc+lkLy1Ag3yxSWcjb1hj24YSNITcZTiD6sufysechaxio0In
bbqjJySjqr/tpKUpZYECnzQs6gZH5kgZu5NDsBv9SvnSSv2F5BmMngJqZScCB0/G
MFJbR2b+BEOVd/ySov90xsAIKNMwZ7Adz8tbvrWEo7NkjsZSFFEkgeNtnyVJbzpm
ddBc8Sdqqxfqbh1489vI7FAv3H4FhzrAXKQyzYYZ+lGaTD8xMgR8AFdOFRO+zuPy
f9TPjvjA8JWxaAOPFM6IcwXjOQLCKqClYE/TXGFL4adZSWlYIyJzTvFIyn2tc9E8
t7B92hBtdZILib63O8xMiNCSKvTYPd76gnqAqD/lvBi1qgfWWMDDDVKlOCFtKSX2
UOX8m5wVPfMUwhoNIZZG3P2QeJG7riwU83822+JJoHx1ZXbJ8L+w7472myXY2H4H
EmlmP6CIzdHlSl7o0srSBD7GnbugMszVlxfg4uXkvt2RgdGZmyCqodz+70yHVNfW
sKvs57GXS/CxH29t5JLlrIAxesd7h8/JovMTXORb9TL8/w1MHKNDgFdcghQ6sUT4
iiQMgx02GxUT2Wh/wkDA0Sax1vxkz0WqQQnRVSs66YyrYN1UdHXbHhnyf+aBB56o
cfW8kXf9wjzzBPmgMSdl28zwugmGjwNUWcgGYXhKNCXUuSvGkV4OjAhHE9PkkUhO
ptVZcbMXFXXH3RdwrlR/2mXENfaW2KU8+eTKikHwWC0PK+HH/ebvgry3zteZgPD4
PBi6nSUx51G88/xbFi/jo1s5M6QUfwVb4sMqddGdAl6KnLbSOrnVxN249wFTJ9QI
LtmV/NWSwlUDHNZ2zyp9M645foJT0zWM7aWfD/rLGQggEu2V25ftVuxfz+YQ64c5
ol/9+IglZw/QFq2qmtFusrO+aUzDD/G73Y/bpl7KiOQfz61y6kB5A4YLOBRzI4e8
t2izB4+rDhke+hh9257yWwCFzcHqCvdKKsDK1adRDHkKwb9W8vByytvvsDDSpSjM
YkgcsZqp8ACTAuDljb4Jt+hQho7WuA9OVuxBdc6RqJ4VrAZ/LensiwiPkAzHkG6W
Eo1InqNXyvM9XfsqS9BmXvB2n+SRzH2aswGslQ4rq3Y4WKJffCDYamAM1TNNj0Wo
RxRC16EtoZDWVKmcHvW15J6SbmepGd62Rbysn2cXnOxi+p/lnvyk6BvCa22KAKJd
rSbJK58LzGJvZ3pX64IKPZ/Tc6c2doWROs1i7H2bfeefZ3GmxGRlMInEOnhkK8L0
qR6yxk8E/1R1h8109Z9WdipWmAI6P4BtYTC1MlEovgkXSu+6nvvcBiHHTHF87o1N
qjNUXsAt91eQmBvlUrH4jt1KrpGcWr8JqmlurLn7x1uD6uwIIBtIyRqyADrVXv4i
cQLnfODzsmtH14oFWGEQHS0EEMeenSP78ZcDbnRcBXdzEyR9b9d+h0wPzgcQ3Jg7
oboOTLBk7fim/tbyJ7JWceX5xrFQCifPT/cYjSreb5CzyjjElGZa4tIrXJ68KrYu
OW1WmSVPilW1NhWRUBsZiLRbWXvPbwqQVw8wR3cKq5pyZjgAg7rwVKE1nNU7Eni1
7X2A4pivJT+Xw/DK5FYjpu409V6aYW/O8WMPkyYDQNwpZ2tc/1BFmOcy9K+lp5IA
CT/L7DrCS9ig78cZgGpl52SB13LA39+/Z8he+jFXrK3M513uBwHSHHiQgRkV854m
IlV4w+hmo4+lbu9v++IUBEBC+ux1MoqjlDZ1byM/zdIV1iXIBGChOQ8yLMYagXzR
kFVdh+8V2eFQw2qcBJ1oAlk5NjmQWd8b2Aj+IxaXoxKfrOQGCf7pVF5S1byB2y55
ofReJ/8mH4gQh/LEeBHcEP9aXzanPfEgaCSo1c0tZHuEugV//E6Z5bNPk6JJKdk/
s24UjbODEjpq1zMoaMzrSyy2PZshBMxi9r6rCnYe4vjErfcQsEDx7ohrx3m2QAdj
R4fhj3Fym04Gw0ByhCKwqyPqlUMruUYekT8zkjjQ3iGI6CBhKSWtDfNEILyryHUC
3atC1uwuIwhUKEA816VQhbpHrN9LXbxLZXE5e0SYswXND63CdKu60xLxNmOwOiSg
jrpi+mi/wf+7xo1Mu4ThyluyLd73i0mfPo8FM2WXplETYDGO/mfDGwag+S9/Z44O
tfwXjD7gPUEoaTJmq4OOkVpJKTBhDjEcOBTs9dVxablfgd0KOgrmmMV6rCGxZsZd
aoHPZlcBHWNC5JckrPbmRQQsteVgiMYriJ5s/EfhSJHhpexuowZlhnTUS/hU/iRk
QaIiBcKLM3PRwBi/bwPOrsg7+xk6B+PEJ0EXGdleMnbosgV0SCQ9N/E0iz6F99To
SknWJSreWTBPuA0c21s+QFyQG11bYMqG0rxv11pBcZESMye1PwX8CRA6GK2MTZa8
fbTxO/PKUF0/UYqQc9slcH7uH+Q+hiLRUTlP/5H0VNK2YJFW7y0fvFP8LKynrL0Q
jS//Sb0N1uDQt8rcM7xEjUbVfX7jh3v9x9sd7tV5spxqRUsTJkqhG0xTo0dcclge
vXTX3lBm8giFeLuUpkN/ZrFWe3zFwvyvie25cozw9vbjDVZEMaG/DBd1c+w2otIr
GBuO3A4/u/KK6Rgcd6MWJdNPFYD0QTfGJFjwefRdg2YtLJ2Me4pIaoLOboVq8BaH
tLjj5JadQTSBGHiAPhWRA9AvFb1+f9EZy5DKK4xR+39sesa4BQZLuQYxsiiI6GIC
9k7lK9R53ThUd1NbfciFBOIJv6aTKYk5L/KdTNlo7tadUJ0LppYJs47NfYgOK/dE
W1NR13FYTAD98u4N85Qu3upka25zL5nwNIq4z503neqzw9lWCsm23v+SzeyJtH3/
ZuR1eyTofxMX0T6sTUeWJw+pH6aywRIWcRI7D797Yj+y9l8UY7ArLnNHFY94EsEk
YyWaEnu01u70qsnG7UFhihz/l3XAWf7XqgKdldMol2vr+5E90CTtI+5RFhEX8Tcr
KnYC4pzb9xgwrtlwFlNSxDyiX7luDb0mEwFWtXH8fM+jL2BP0kYeMNWz9crkyybL
Q9nDShwXEmSHWVA3i+hhloVjyp50sjjIptL7lPMkbZcw8QoFVURGhhoS21+2My0Q
A7nVEHf2HWkhHGKOoMS1J/IcEvQijuhAQxMVnsu6j4AxnsCo99sqXCyLtmgUxXGg
GnD+ThYS/3DptkYGWxYtJYJihHbniU33xATQ0Aj2b3UyGjf7fnPKsbYo3ZtFX+58
ZPWEPXTvBXQX6xzFRYLvqyJLm4QEu7CACVp/hxQ8Ojw9lcjoW/coCEPmvZFwq0Ee
R/faA7/TGXg+27CByEJakFHgFut2RkVmJWVcrl0StUym3soatbfsB3YXiLfvW3o3
aKcYLtrGtIUd96KyndL/XuFN5UMPnLhrtq/n9eIG2l3SBaIKEcRep+sTQPKJhP9W
CqMRoNEF/Wk8BbuHC5zGJ6T4C7CPaQRUNvEGCrq5hLOwLwdkpkAaamtAXB2Njg9P
OsnEHL+RaQ+CQ9vic7bu9RPQi3AsY1SckhndB6C0b1lhCor+hexTgV51SVErVO4d
BUxvILoe5YACdl1HhXfLgiGj8j2Bma2YO5Sfu21h5ib+UANwlynpu9sV/Vi6wL8K
Q21B+zFCjSE3V9Mnnk7RQpLadrn9rqMwnM9sLQoWWFYnWPYPwTTJRtQ3S4vJJU5k
iUk8Hxfr5v55HogaR3i+Jp6fH2hpkugBT3+xbSvo8hlozn56gF086OCBS/k/pUH9
hTId6GoNAHPRHNVAX7Vpw0UkkQHz6gSDFYgiFNTLNaHpENSIomGBt1Jr26KNDOQS
KBoKovguelA8AFK1laB3YbD2RewrCNow5ROmPtt+dWtEVd38hP20hd1g4yv0EJV6
YcHO8pslwSEor0BN2GHYebZtMCViGpsINnVPaZFcnZVnXQYPvW0ZHU9z1nrtt+38
yLpePSQP6Fx80XvojV21+Qk3OKCqstgato7dLzbwAR65V+WmpDR78FMCZkm06IT/
kqEifB6LsJUW5YZ11FyXuIhYWH7j+85lPLqp5+uOMKZggj92sf4vc9LsidJpN1nt
+s8qB3Xzc4WEvQkWIYeWp9iN0rMapAsoslRcCQDvJYCVjVyIIEqHI5gRev/iPpdM
qzrTDu/RnrK3Gz7ZHtLgmauvY6a+iP/xe1tTACuuUa0ipyDj4KueQsDwSA6WqbJO
ze2AsIRBkvMT55GH6CsRt2rNMLaiF0M2ikrOeTJBFfrtT95tiid4HVomftGNsWFG
N5FP7/gDl+W55HBr9pn+End/cSMmjmPJTu9nwB4wmzjEok0I+AzL3YAarN7+KJmF
2I+YqHH3EhJe6cUt1VcGyeVBZa1BH82j88xNKni/CwGxhtLAAVJQWLnZnSoX2LMW
AU7JYD69iSk5dS/3pHaiDtOjwsdlrW6V9PoI6E358PH4tbolHEYXGcCUvXJuvBTw
/XvYwX2K1IrjxG+PvXbUmaOCzdi+WkyUJbQXlza9P1BcJQBZivY3EHaC04JZMRIh
QblBB/jb4g3hhZ4t2oy33cswvrSWZNovsNa8Zn4b9HbaEy7kSAFLXrMZzEHcuHk3
x5uKMnR/OJxqkD0PFCdhXGP/M/mg/Q5mWR9bV3ArdkxYuvuyLx6z41p7ZuA5SOpj
loyP677/amOBO4Q87OOSlj4NfbHAaxbdybXr8xOOQLhEWtac4zeyhC62K+mpCSaR
XyzZuMTBNIeH7QIXOT8fi3fhLPPHUmtEhzZerYGyZno4MsSYfo6d050ZS6kV4N/+
fPqnnYk1j/JdOy9AjAu7OXSaUeNnD4CMTbfy4PYZLF/ymAYwIeLpYrBf5IhIb9dY
1f21tVpF9QTTfEzwLlMC7yf+8DTjl7b+QlV2s4pq4GIOfqllmaz4h+4vtcygk1Pk
w60EQqDtV6gb4CoKPXS9E+DmMqeLeBs6tqbNoCOhEVgH88O3uiOSSlXMlqwVevRx
EGQLmrJUWULRJ5v4RNTX8EarT231+NPEQiq+nomT04ALiJsOOEENmIXntRLUoOEG
Jt1FhkTk4Aw7DP6Gv22bAKryCEWyFMGsGjjo4u/cCI3qrUiHdYneU8rv2rtaoq2X
lUX5wqqyvjg9McfDwywdbxhMmUz1n/oL1A2o+7ARJmIvQ1zBJ0Q1FnRolt03OSmP
zASItnhfFcbgXQKpMce/tdW+ASwRpeCQVlXQrMB3ZYXyHDHpB50t5YBP4dzZ0l5P
/a2R4qjuS6vVTc+4u02vq23kpVFT+5vSPWdS8CnRlwXaTKvmTf0PMkOnDf7oMc1/
SLSnD0xRx4TNXis9ouVtag59yCbClubyDykhnccPyOSzlh1SKKkxtwymsl68Pzmh
NTjOnN9J7H4xkITQ+iBEGhucHBmrSJkHqSmcUCDtq9gyE151LAOijgd8mvnbAhJH
KWT0UiOWEyC/Pm4JtiGlTr9RfzRn3rqzvxH9TCoN4asSS+vUg49bEuZgLJwp1j2o
jcsCmihJqecRZS3xOGbgRANGR8/hAb6I35DrW4b8cv7r9HH3xUKNi2jsW8BLQoGa
l261u3DALCyUa5vyqn8HszOicI/S3O0X1DTrZ9grNhCgoPHceqW+bYdo6LZreChb
b4q/fJpUtj897jcUTeOvlVUEYQJQiKmRMSenAVkcwc9E2AUD969hYAW/WxId0hHk
tBvGmF9s79A9edD1k7qecJlvrkXgKOmwExV1XmOkbqAFmBh5VP82bHy5t/hwMev1
uld0H0/2XYoLN4la00rYHktdj9r7ma7pV/1/+GmqmXL0H52Ye368TGd6C/4dODQb
/QLV+xFmMap7z+wYHUYXHzfZX+f9tN6mDqXT8NhBvgxHLYRkGg7rCCJq8QVN3wZk
dj7etH2ALsOyVR7IBpmxiHg3TtpN4WCRd9xgRpCIrhQMpos1dVCdgu8UbVSdIKBy
QEbB52jwpXLuVZt/SWSiWzhtg7dLYpeJ0sFS2BE3e/svpboVcaq1mEJsiknG0r6/
byH1QV7cQU7mdl75aN6nRBolxtrJG8K0XYhI+129be4WaS8Owd8lIayYoaIhg2as
us1beb03e+2a/MLZTuqeF+o55xPVRnU5XOtoGKi+2U9etEqfDl7VCKr6CF3959N4
/kwZahhXaGTCo/56wWHNtJWFwUea6BZ+mpflDcMgX+wYgBLl7b1c31xTYNjlSjRr
B0OGxiFKlOB/kd/NSiXNkucMy6bD75I2D8yKS1J9sBdeFkITTffU/qpyaiwRQmhK
eDT1coyxRQB01R6FWAp84h3XigSfuI0yqDH5QWurwsucheFdPXXbC7UIl/BcamkU
zzmhNFUFNuXF/8vQd1GvSzcSEMisMOeGnfM9Mge+BWj0od3KX7ZBUQ9l95J2e7yI
g2BBCsSbRrCtZ4wqTlDe1OwaVoxU/1MPtJWKTH1wdFq/Mlai2JIUcsZazJeQIUk+
8QJyKdRd2oY/RVNSmhP8BbBKLiz1OZNrFoC2NGoK90t03dYikYJaEoPQAaiQQKde
mHN8PdEYlXnSaAKm2Iy7fZRg9NOZp+XpFeRow02pcnVrSpdydzq2NVt78lFVHkPS
KystfLeH4Pltl16RSOUfiY3amipz6MYL8xEJpkHDYR3w00Oe+xbHPZ3CGsPf2OMQ
Ip1eSY6AkivsPsvW77CTVDSJY/rmxEXldXHdpK0rDceB2b5c9jxN3GhKY7V9tPTS
MpA9Z0Xu2yqE0SQsVSQmjQMGfnKUksRb80toGhTvK6mUuZWgkkfuqF4lWVHrgF4v
evaIQktYjioSa+RolwUHhKTIuh7E+AoXc8VSW9OWuObYQUkJgbZ1KUmmLPMIWF2u
Pv+wmJ9LaajhZAmX8c6hp64qVd6b4LZ8Mg6CGSZ+Sy5DEaCkX9+Pi/V/abIx2Awm
68VDFL6Xm2iVKse8deRbQLBF4r7gJM+QnjqQEw0KzisDAseCmbHl7nNuDNYuAvrh
TlYFKQS6nIV/QBoMBIfoeOOEqcLK+40Uq+KsqU0KarFDtTIqf4VLVtMRBmqTmbO8
JxNfRXBPnDF/bLYjP43wCeLVDxJJABuUF+esGnHxjrViSNrmGTheHit134vRTkVI
ymvDJzuSQVEMxWzy8pudssnCzrtO5rWDcHggZE7xXHfLR5LQ4BIU9Keg7KyGEq7U
fXKbi6m8N7VhFGy7URYxwpJneiMKVjMz7ESvr381g5XrKSUbRPMJEti+Qooqosf0
C5gsfB3OHYqLVrisVQJICRJwwmZDwuI1VvLASlG8e74os7toR0cdBbTmOw9B5dy8
xjBdprMqaVIAvVIP1ROoyn4DGkZEYxHMf5XH2m/hkIjrGTlmNyrcmGCKrHl+Bj1l
KU5ILOFlMpZGY9/SZHsKI5EcztPUPBYQ/Chuj1Pd1zj9QKylloXlMTvmDMIoqIXu
BVMMrG+6YtHNCZHwuHR7jSjw0DOAwAug+6FktdwK2CYkwK5QWD1N1A1pozyZU8if
iF6zW9+eBSc6FuNq9eXj5GYm2pN6a3gx8mVype+bRvSw1s3gE2vyzDnL5CTAp67g
4XCVN8QZ3lnJQbfmAPXzeD3N92kcNznWrNFrElCf+2yRAxwGfGmjRpbm06XobDkn
+GXxkVzTHWgVGxM7f58nbHu+Nv8Qi7EaRA0qn84yyXvx9KJmczjqP+TvkduYwx6t
K5LuttMYu6SEorP9eVo4MIb23PuKdXLuMygobWOClolz7sjU2E6SI8KWA4btRBwb
MFACSQjOTpQgwO+iM+uvksJ5gbEBKcFx+Sulb/wdwPV0DDmhCq653XqeiCn9xWT7
KAHixx3TLlqfdTwZ4Dte0AeOK/X82V1jPBG/FaxOCVDDg/KmXj0IkNI/w3nhRPvn
xXLHnQUa7gCQ2EVk6NOtzGmjewYnX8tYaSc/iQwAq6qd2i612AnGlN997hJZvWZf
abHBUC7S/T1t4pkr+XCOvLzF1YsfQnxtDEz1intE7vh8iyAAkq1cg1o7XDIXztGr
5q3N/UuP9qAV8wZDyV+LROt4ldFc82vNVTb5mz1K6uzKBUgAM7pcDYijXigE1j0f
KyLr0Jh/MUAdpTV0oAS2JnlXmraqBWWzdUuifCgz1xsHtjLF6CYYFM+XQImR9vgF
+PDZwiPLMQMbirQx+nFqacJ3KRTVqIRqywXB3Xv5JBDTrbD+HQr2fOeTr+vnc6Xx
iRoJrRrXRwSLm8uoEc5QGhg8BBFJIbp9NAzIQy92KGVEurBliF5Sp3k9sNEBYmul
E14KcOYaMMF0UnGywNld2O8+HiBnBe2w75opjCiSkbQGFgU3qDzfbwzGRjSGrn/h
sbPiWNmBJXwj8GjXQfIoqpuHTaasFEaHCoTTjcYlYy5XCpWt7Cq/vFTc1ha6g4a0
VF/JCBSSfU029LyvoaVxoXh6o48OtqT5G00qxS5Jm1nr6WiQNNmycE3ZSyWKlsih
0Eo09WXcbxPYrwfnQdSAI/bFvXdYs9o7ruvsUOsqu6lh5XdWOn3jFtNU/HKj4i3F
Y7tj+VcLXwlVuAmt742CkUNx33ylDyuTojg0w3dkLEPmojpgS5iXkCmCys771E4w
ExOeZJQNu+tyvPgu9PbrYl24P8nd2IwakJmB+9VF0CNYcckhweVaVB7kjudqpAsO
RKHGc7ucFRHBBfwyOC1ypsp6lxtiypN5OenUfVOCupHlR/4SqL5RTKRn6QMtVtYF
3nZWLeULCi0sP/Yl89Hk4nuc82JXjMNHizaqQ4QEosOAVudhsT8ZEqROlH5NGogQ
LQAjVtnkpYSJS8NC+Y1yymOrFYIpj/dKvdDXkbSDELe5nd/x3Gg1PgfHrrfm7SAS
YBAUM6ZTzDdBN4XBA7Hoxjhi+9S+JFS8QC08opSF1SyMiAHQ18VEWhLGluFytlWS
reyZC5LnBYwA8ed3+mcOTSSH7Ojx/7uypRY9EXtFeU6OACZUQdzVEM56iUkFMU+j
jKhUo6R8SfyVMqOwb873LHVizRmUXjjbzG4jILUhfOsi1bBxd/1QsOf7RNLrNPhU
7LGra3GBJ5QCHKofAdzVRKZ3NfMwmJWIwzJrDpDABNur4WE71fTjkuxkJbn50LTx
jYnuEd/OsgTjD2l+rnLz0ml6a07mDI8wWG02Jy2w4OKnMfjGyK7BCHx8XbAwmBwF
yn5BJot/8dOP2zj0/69MOwHpfZo+yNHIj3vKBrFoYBPEcsSP6ctvGmHtVAb0KISI
G9D3Ccs1VrqC0dPd38IfeGnacDHjKvGoh55xobFgtpnO4ai8j8VsA+mlNGguEEuD
uOPjavqHsvx4/hJ/GKYV6SHoIMy2v8ZaW4xVGyyYezAg0evj6aLgOsfAWBuwgMna
RTJ3z8+iZqEJzb6qYzDHx7rn9fhCvXyPyOeESiCSBSWH/7TCsrkA90dTBpN2HuiM
vlIvc0fW1/U3MmKXHlTEcr47OsptBuQApR0/SfgoTWzjSFDFqhAkvSVCVA5f5cP5
LPRx4NqNblyVHhVeESzQOIUTPI33eYN+qoOidrjho7hhcINdl7Oy3d32/tCFjKCr
2Qv+cLnxizO0lc7yMmotdcJafb+hCh6g2wYdoLGlnVZybphOLL+rkES8lsblJCNN
3cYHSYJPIodl3QoRmyjffaKmOZ3qBHafiBvJU8Z+5vSIwmeEcmIWqNBOn86UU2jW
RBfFy0P4ZpIgj0dFjnlyjOE6lorc+eIKD6LWQRUuvwTPZIXQSmFcNfG7RJDC4UUW
J1xyJBFsNR9S7Jc92GY36GxKEb1p6N1CflrirRc/x9LVlXv63RNw5J3NQ+44fsWc
rj3Q+sCEzujJDY3YIewsmi08rAqriUQKedswvRa1z0+u9DoVu6ZnZQQUv1T0TCwY
hY9cA1vJe7BIJRJih1B1SmgwOE4KS8dFmq6qzsJjUefVIAaGugW9XlGQZAIN5JzD
3WZa25z4HR1SThPdz9Dl0bs+4zLAYMohbSJYSVvkViqMvu2wDxCH9Xy5YQyozC+F
xZut1EmrQ7WTku5cHasjYSsuWckOP40oGOMK39R+Ydk47uo1Ky3Ml5I/HVeTSYsW
gwKfKezMBZkzmr90FMXW4e7SbgBXED04JQct3ZjStftLNsvoBUykv/xnWJsS5fZL
mG++YJQSByMpYtdescNCyGfDuZyggdRLEo0c6LPbfRmC3hdWevJaU59eFwJjzUZ0
A+99HHU8Jq1YZW//v+/E6Vedxe83fQrjkplRntwJuqL3R7MfGWgOSRAI0KmXneID
VPjhHT8dxOX12Azw90LAbONqD17K8bM7u1z3R2aCxT6ivD6hNj8sQQPv0Mp9LJ4p
yN1QUuHtExXb/MiCJmbhbp+fTuFQ58bKXXHq1zc8DhN98q1AJbTTZe/+5CTZSIw4
eTNhs4SyMm85fAEGTsbAdXUFvvhc3U0h+8ThbtGo/C8NvlEkoo4wk8ZrHp4Itz83
i23hVWEsitMPUHMww5uMdmUvf2xm0i9hIQCjjuGJMnKtmPAjB6vDhzdLolq8t1Sh
SFpchLPf9eITtIw2qBqME5rq/St8cA+L2O4+2Yw+9Bn8Y4G+KD7khsDt3usBSLcz
GAoUgNvgd+zAR78JwSr7LYWyGhL75OrW5QkZq1sB2M09Eqa9CMKqIz+z7qFGkYZB
MiZqgkUi6EAvrx8Qje8EtFUzICZ2bxajUeQxxRYRxwBVaJscTYwnwjInSNd/XSxg
83DjYp37dbG77OhlZanOB6eQneCwdAo376Bu3UUhv3ow+knVs7BMTnB1tdDmjJVB
hIKBqVzHVgRC3ViND2VFujsPancmXk8mirZ+vG/2n6jwVFF9Q0FdfvmEddL4pphL
awtrNjN0dolYV78+wvHaoquT2HeSvKueRh8t6/c/+VLF1bMHAPe8ire3dJ+jh+9K
n4b/fmS08W7cp9GUa7UPEFZuJ2bYQI+C7AruzvruOH1SvisTWEX5YBouja7V1XCO
qsdWFuMeWsxk/CIFYn5ruwLuJSNpo0rkaQkJeHhqUNhJGeX3FOGksKouflJ2Q+/S
eT4RUJcaoDaQJkMSA2F3HANTiIelqK7FJLe6bOTAGfqsneFOqhmyUKFZavk9YvZZ
P5zfuo4bYXlK7kmC64iPeFsyNOA57Ej1p2wB4z2MDeNaCx6Hzdd6z/X3UzmEMcj0
Fduqt3fGbubSJ4hvgHW/48nNAi7I97ZOZGkygBNhw61aprflaE11uMVQJiahH8/b
tgzcdYAqTcFWFBlc6fED5M74OABVkGBGnuQa/28GaCAiZOACyBMkdE7mhWQiG24z
WtcwbDwt+l96g0XpZ4U7yCQnIcbBRxL3mUSnQNwrTriIejj9hW2tFWKvwSTiFYst
ypt2ABjAXmTtvuWiAiRNfbKEb012+OS+KAUHBVdD4ECYAsA6jbQ+Z0WNttWESfah
urr4vSq87Up5hKlGIGtxzJwf6JVjoB+wi7ndl0aaleraxR80N8bcctLroU4FgPGf
orIGbBIebPoLFbU25K/9V+MxydMyzpP74yksnDf0g/eawV9auZ+0cnFictbtTxbL
/CTnMmIh8SnEqlRp9Oq/9BsXeT0fTQW774qOSmB6+r0ZMDuYv4J8HHiKDyDRhpJR
MggbaljgN8INZczBAboniMs1i0eW9vVc5HzYjTuuG7ZffwMikyXowlKfeMWk8NoN
Cq2dQRRv/djTkcc5bprRp6N9YYDp/OQcK8I63/FKY4W1KdaXAFoC5pLq5BM17eYD
VgOJWtIuJzDJDlWK5pNgjg==
//pragma protect end_data_block
//pragma protect digest_block
XESoq58O5+8tD2kTlxdLBnzTS7c=
//pragma protect end_digest_block
//pragma protect end_protected
