// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
t/448GPxsZQlb+zCpZshtISJW/mpdNFghIffNr6bzKf7q6u4Z2fjN4l2mHlVPyTC
9Br54GA8s8S6Gx//EUBbmLmf3z12t3PpV8Knf92XPSjTOqeLZri10fqybsVaJjbO
7B+kM5BNyRSKDr9qTDh6fc994oIJwa80cgs3r8KRY+ArBeYIbleB6g==
//pragma protect end_key_block
//pragma protect digest_block
3NdrBIkihDrUWjTcJa8Q6v0+7bI=
//pragma protect end_digest_block
//pragma protect data_block
RQy8rgFJb/qKAdmqxQloLS56kj9M7j5IAlJAdbekZYadJjh9xHUBHKFlpzuW7xDw
1u1ge06jyAgUKg6rrQ75wcM/iYN9vOhAqBBJDuU9BZdq8OafLCUG+cppJAsIyBdL
99A56b/+ZooMv7a20+wO6xokndX8YnmBXAnkYcWp4b+pA4X8GKWEKdPWLrU/Se7k
QH91eQ1eGU4H31rxckD/U4uE6cy5yFsEZ6wzW65tBsbE+SiprAud9JzXfkV+ekBI
piciBtFguiM9B5paJFHmZraMaZV6KYDj5LjTWd0szWjgX4D2NLpuSMdHGg/NcoDF
iTgDE+mQ4VhUMGaUsn4MlT34J6RYBtaG+5suX+iElpdlA+er1KXlu3QsbqtfZEfe
hbzjitj+++EuyFzb9CKqW0hLgWIUzuyCCjNgYAusoGT7IPAsDZAjIcCSv3bjnOzA
0CQCRZx9Cpu6RQysm6rTwtDnjYLF/QdLP0qyWYLmphgFc958YYTBXhLnlAZzp4mc
g37T1ujlQUU3+lqEGci8NsftTxktriiCupovqSkGLrpm1xp7r7VL9IIQCepre+uQ
2JI/2Fh9f1XPrtvPZRKGZpkXNruldXBPgjCTpYxadaglEQWMejMKh/8eNKoeH/in
KdjvB6ljILnPBs7ifR7S8DzPpp73suRMqbWvYN0VijUvC0wDw2eFWyYQQSEpUb9N
WBzwFWSsEr43y60xAidywydd1fxHNp7xJ0xpi3xi670m1gZKe+TlaWdtr+oQW2Gf
iViTGEfaWT/xPpplyggo+E4S+sxvmPwHjNqBPAN/sofUvH8A3GY3dR+RJYjAsdq/
FPPT8CoD2O3IxXmSSgwJTRSg5kEP7RsxpwuPgOp+I2HvfPVZquSfRQApK7sRleWD
mr6hLT/df37eDNE6DaPIZCA4zKEMoAhqOHk/kL+XcBVgp+WiGR3cOc9sKa2nnRyR
n2a8veQGunhhUgBY1PFwOd85Sy+/Wku9uSARXmtqcw3PRdQUj9IiHkHwDuKBVryp
58lasCTkvEhCVngf0zumBO5YtEgSHSMwlXizjRGwg64SQVGXELubfFCKkd7ICFoz
4X66pCl/nlM99xswKWS5MbpDoMB72EnjimgRjoKmTYO/ByBAWadehGTi+PuYAHqK
zredVESkEEapax87lYpSlTI+dUVVH9SO23AmeYXANLszSR8E1Qh6+8He/P2zhPg0
gs2DUmUb4TLrWuYj1zrSlPgQZELQBoWjKrMHfmRtxuqhJ+l8rh8BGBsgYRmAcztE
0GbR5b2Fb4FQqVTaWXiAeX0ks7SUx5RdfBMJzuW72/GXyYCvjxV+2a4RDRtnMq+E
deHOgiFfsOjK1H4/1uS/wGlfTgGB0wSyQ3vNIn6ksD1mttBLNwkwOe3RJCDYnVt6
vCSlWrF5EI3MG/UVySvpXJcUDKxONzqZr+LAx0H2vu31qV/20hRYOaN/av+uE+cO
W6kdIbvIB+Kl6+V9rLO6DRWMagEQabw6gdyI8wNqv6jB00BgvmMVzKfKTSB52Ftr
O5Ze1dTpTXLFh5d4IBbl1GVFk82+XJcIAyoflwXfJLYSzaHP40ro9mBDC4uoJOUu
GFbn3GqWgTcNgkBpsrLJSlmTaa+4YTzojd8PqofHUT0qaf0zelB0v3dZSGrzhAkq
qhT1/MEYyDdDVbOP1oA05JS5U2vmZl/wHLw50eJKMoQXnnGc9u83UoSgBKfuAoBC
F22O/zChuMn2XifCs5qPQEUquWU98uXm5doG0f9xLjm/PeNmS+bSBWGeEAjlOdOY
vRtHtO6PZTEEe9iMX0qmYSLm+UmZDdCFT834n53LbeQYD5Yyyzi1AgSfwhXETiRC
nhHRcogCyTkfNDTmF2tWriJwa3XxRVUl53Csnc7gsHGCP67T+QRT5L+GF2SwYhsk
oqY0Zznz8YOmVn98PTqbrObKeDhcBHiaqS20h7NtifSnjh3mA5GqNTN9k/cecwjk
y+4SX9BPQ0hpqWcUjfZ2ycSGGqsfLQsquk+03qqp7wilWlE02RYEGot6lVd7gT2I
bRq2AM4tocxnvH+fEuis9EcenvFPJZNUBcbI4ZL07L47736w23uvftAPb0p1F2hQ
eW4dC7dMEDMJtZApmAPqPiMRaQ9vGxUSSZ8PcfQ1ZC9kWhiPm/fjw7UAHolAusAT
ST1VEOsaB6/HpM0UTb+3NeghWWpuxZpG79Tn7M0m9swM3Ig+sRbkAJfVyu5rabNt
JDzBOVYEsBfuXhCX+lr427igOSHDwgLjfaHAkk8k7C7IpiF7IgbqjZXHJA2GDeY7
mJX3elw5qxdrZAt90Sv8E22D2a97bpfEtMpw9Gwh1WAEn89OoBSQD2+EsYbIfxxT
GqJIpxJ8Vph6TYEjqgoeiXkUy3VKBk32iBoSxVuxjoJBfG4T3FcI10tBxq1yEvW6
QbIspJkOtmWj3v1Z18aU7H2uqjnH2PL7+noPp7eWOrZzLvtY1FDv1u5fnarJV14F
NsnM7tQlUarCBVzYsDEFD56RBelzW3bAsYyCQKSW/D9hDdRDBc1h5ibbaxsPa3pa
BVaHExU8gEYZTgrB+iker9oOxLU5oGG1Ed+wwfk1EaZaNjF9iBR8cNwjZndPUi9s
LXWEyhWaFxUbu8li1aEHaZRVerNoesFSU4u49lJqhRbf7EgjT9L9740Vet1LL7m9
uS3LUvEpp7u1IXkH9CNcJGQ6Ehxf4d5nyQLx0cMt2AquMMhLF+wbgKTv80Jp1hnQ
CWcvDQYcB3Ki4kl29F1HVeHnf76IqdSxjR4fa0LXy/98MyTdYGmbLpEAKlJ/K1VV
NuuR0eClhAaJWrOqtIktF+LePNyj01qnZiTPrg3irZ/UT+5kGauwT3XAijYLkLxh
CNsIOKgSgbRFLq2e6ldg0dP9k3XeKKjjOKW1qq18XrNwmmmt3ZEQAyjd+13JAQYX
3plpZZQFGAF5I6UlutcUE1hYgNpz+uE7qtOjLNRlW4utqltvYYlptPmNqwalyUfT
MQGEih7XT8hG54nZpqxW0G2mKBMnUWi0eMZr50T0ytnbDw8k93nf9szvy4yCxN13
7tRJ1P/KWm9uy724repj8zeZdw8RYGBd6ckWm4QrrRvuJkl+S3bgh9UrkBrepslq
djGMHbYSqSmVN8i0RHZ8VRZOkigzevx6H/0F0ewPgl2sFD6Bm/mXM3U6kiykiM7g
YAV53IABWuBvqvx9G8vNTna62Z2hAzmljjduwYC1lqXaSVrunGQifgjp7Bge/JyS
gAoA4u9zicvpI3duRyLz9BLQ/U38cHPiG7UGjbPkXGQ3KzCrZtDp207VyQUrOSYh
58TqUiOsjymUeEsB6iFX7xv4edPNGoFwgkk+JPxQUUAOL51ezCJSPKoP93XF4hCs
Skr0HWEHX1LpCrobkm0WJRlAt+myU8Rxl1b2uDRuvMJSnIEtKNJEbuU9zXlND4BP
jX2usWU2GlU1nmpWmLozkzEZrKildsqnOCENSaLSTi29zQrHsDB/lV2zVGwxe52B
+QAoiyZlf9IxJ9FUV+S01gj5yHrxjzY372bNX52hmdq0oTByVMmXwOpnURi54MR0
SIFxjJJLPMpNyej3Sbb3/BHlX1/NdhPptVSMvyKt3GWR5bpr5J9/+f1HkHOjATKm
4h5KrFALr8wchED4GCLLKlVzv25LGUBIYsmc39NdF0YaSkVTqoi/4XqtRsog+mgV
IAUMegKxt9cDojmjk8T5jeXIEjQSqd46nU+7ye2uShreZu7c1Z4DrJolIUgOKPVu
39SFV+YFER8F3VtMLAoHOaxx0Yr2tPxWLa1UMqxCjaJTxvuO1DwSfzaDaPLIJzu3
Z23R6f/w/uXlr6/DDw3Ki5OvxoLGG1xoBoAjcHHKxdu640FlV+DZUJU1gbAQmwb4
1EFxTY0J/NYjpJlfMCFTJ7wcY1nqBjHl3SicVtn1m9TWyPtbGFodkg7EPcBkftwU
1s/neNGI/bqw4KtV1TTTKm/sqT/nIhIBvTT4QXze6tCqMJXbtmFnKoyrVCYALmGJ
tzPpohlfXmf3YsGcc3pruBgpLN0WUQ1AHOxHvgXU/zeVOyoyICalcsBYT47wntz8
XSOQtrphzTbZD+emfGa86Agz2y1xxUONAwgqpHtwFj6rjvOwoXdX3VGnxEBbdFXy
2hRZGp2M3ap4GNXeZ+5uR/aCZgPcdH3OvNaYRh5ZsbPjMuBPQOTjZV4WdWu1xUuk
FCglUBriYPQ46XHoq3nOm2ZIGgKcE9ywhEkKbni2n6hktHq7/5s8g7WEpAcJZwuu
KMwC11EBVqDgZjgwQHGVV2g5Juj3FAWsnHCotFTjGrfH+KZ8Rr+A5KMKEsMBAyWE
LWdWkidw2GKBJYzbv9jr2uXwRcOL8hVLrBoG9e3UyfjoSpj6lweTkD31axliEnD9
aUmwkoDFakb3g1ejAxbscftgNvSq0bHuPsgyomUKEYAlhCc1IVbrHgJRojh1IpTw
mqNi42e8JEMlmJoTS7CN6lHqpatoyARdjIUXKV/70yMrzjZsOG/pE0+xDpY3QmcK
dfSwOMlU0HZTgBNyb3YO6kQWX3E3PwVNaI5ABLmEug6uSFMk+MDlq3RZSAtVqPCB
ka0t+liFFg2eJsP8KnTRJAdolyohCAQ+L8iRg+b/OiaFYRecX509u17vbVpbtf4g
+/ekbC1xH2WX0r8JDfpZNZV6/JJ0F7zEriWOJs+J40QjZzrWfzVilR5NADZr9Sks
IAuhM2HhIxFd6d2BqjXWLCL84CyHTn2veXcgI9nUKzRaqUjjhAOcJZz7vs05RAcr
yOsCaqtWMoYAMnl9YT9RhN6z75yLh919rCp9bRD2GQEYhqS2PzlDcBoIAPxkVXrK
OlwlagUl0PF0A+6t2QP7CIPRlyJ/yfActzsJLgbzvrEM6MuGoZEGy2Y5c12zk+0z
O2zcmsHQ6if9C/Z8jDSDN5yxQx+ib7Fxyl5w0gR2X32AzmU5Tn4EGFTqVjGVSAWb
KazMESNdYQ19hvkOniZHCbZaTUJFaDMaZbNBQuUXrQxMGkLk+PFK4Pfs/oo8z4ly
HPukgO7oBsNN/nJ/mHf7MWT+eCIJH9bvpqF+CPdk/zq2qP6Vs3La/zoaekzGmbMI
4L9Zbh5rOHwbUnDqpmzZCPltgKlgBTU+sZctlGDRgYfNU7EZxhBMPNrm54UifUiy
vMWdjWKNIDYgY8QRDQHkMDwMyLjQrEMe0S6RBbu30xTiQHF2b8jQTc2lqGwIfqD4
45ZjV7Mm9GF/+UBBUeQ6MozIgGXwmqcY/KBBAsQ2hYUwlH9ba5Te4UuzgRy9RMK2
ZoqU5L96CUHUKrUhHgaqVAlS0S0zsxDXxTmWcBrdxaqOTda6ekLD/WOB+LBLYxBq
+DAasUvrNAR4BWqk1Zhk7w8QQMyqtrW73G6WPFsWaSCW7gzm7sDZb/hDDDRHNjz1
AhmFdSkIXZH3KQCJzU7ygngUsYOPF8Ir0uQod5lANw6qTxvoo7EmDo6ceY6wQxhP
EAF9gJiguSyetjEHx6bjZURQi7pd1TEjz/6PP31b71ZTnPjPvXdfjtnoSbbXP5po
r1mXy7cFCyNU4k8uFf2nVkXjB3P+aW3stjqoXLImca7tOk0AR0Hn6oDt7Q0sEQtb
jq75xHFjNgyZWWfDXaPREPj0m+LaHrcwcmCsc1fLD8PGEgQE7C9/MaZ751/U+3di
8w6l2gqjIsoqqFaVw5HmDWjpTgAVFSYlSUw4Tl4OZrsa2XgsOqxUxkQ7DXPR1IKH
1WVSa9jNnFO5KouROXbD9WstYwhTVediX34clnzXaGLTlb7OPybVeXTm5NPV5C94
oSakGbbEt4xv+CJaWWT7CkOBwoe3lGsqAlpT5PeKIb7crmvtN0qjq0TVhSybTxuI
aviwkCCsE+bLJRuEpkSXm0tIvqi7ULau3v0l7Yio6wsAnKq6IQJdmCfOnK5FtbA2
3P/2cBpUQ+m4F5iP4xUdoGVVAccOPbzdiCpDA4Y0XAoRNMg0wN23h/4Jevj9IUp0
goIngMBx8wBTn9k7eZK3VgC21T0PU+QLG1L5nHWMJBVAfsWTq1QmNdg1YQWe8Dx1
f9Er6shgeW+zFnqtbKo3ZlXRZrTKP5TJr2IlMh/26XzoylAcsRjrgYjcdYt2m4Ae
LE3kT9NWk/FiVflLkWi6UvnT2HG50HvVZjWL8pq7exEez+YsAMe8kSbCpnC0tiif
JV1AQQA6WUMin1bEvLRvyywtOcljPvzhneIO13xI5iqnqyMViUKO0jlIpp9BfPnY
qy8Tl0GoiErp06QLDrYBJIuy6DsLgaQMcEqe5l7fKW357Hdxjm0SlcT8rHq6YHdc
nH1p/ZQWcSXI7NMkN24nYF8baIOMw4wp60JfW5g3rY3kVUIXSpcZzInnlxJkRATN
BzsWUEKcj0UGDFRbEzqqrLYFIfQeJr+z4p2dnnwlKlu8CWMzgXrS28/MFVsHSoAg
QVWxr3rh26YVrlrHmOZo4Cy6A6lWBnktk4EOiC4Az+wTge6Bx26kWjZeVqwcXh5v
CjRwoEq1+egoO1+FuzVwXQcyUeNvP8vMU9htxcRPRDmd1hqnMV0ydMoNMGUJdWJv
A7PqC8kxDiM0o9vfWjW89cGWWeVGXHQIoi72jZlEguP9VYHNS41XPtTLXxBgPbpO
uj9lgys7V5QDPfObjSKFgYck662I3bKk9P3+k4a0OvB7ZWXx6KLaJ/ZKo47zFkSu
I1mTrS2RU3Ex/gOW5eHf42exCSOF/CaBpMLVlzqqBwyzYUwU+jR6tT5MwyFGUJ3R
AD/VvVDB3kR9Ci3SSAulnI2vdGawm5LqWg707RwMFH3WeJSxz/MrrihX7Gq8XDNs
s6ftrEyUSGBHRwkKE9PCNSlT66KvtuHUn/elEbiZ6IIxBBHr1ILzB8sNVHeTZA9K
KWBwtxHqGKvKa6oY52XgWEZD+0CLnCAXAFVFe1swNsU6bvXmicNeJhuXfR8c2gcY
WSNTqEZVwfBdbd12mVWF1hxjlTmxc3hqL8YDsVG2Zi9kWxP7V0Co7Am/5acZQwGs
/0FkSgjffvM3nJwJozX6u5TpGGB0aHNTVHs/bGPKG2VYixmxFLcj6rNoRwnHDYMI
ejfboWsAHwPG8JYvS9nRcuvPcg+RwM7E0Y+NSfePVSZ+tVNAQxdLnR1Q1rVbZFrB
CrHcit+5YFIfuAiiGYUOkq+griMIJAloXGNkYUUfNIyMuS22RgMIqmimx+TApU3m
zWFctpNcIoBDJVWRvrIt+SjGfoXSY8xGiFUo72vhjYJR02Abgzhjv+3kPEYzB9gH
XrpdCi3ukwhdZtru/W31KbtVIMfZ8UtBG6ynmcKKdSpOUjb16UBW/v2gF/jDebOd
5GmNDDmQfvYK7814zNzN7HNQzZfRhCl90eJY3l5mERbeSHBOa7HdTWma8o0Wll8o
Acuv1VP+k8/tkx+y12LF3LMU+HXfpSizBd15HzAcCqbg6zVWBxSYXYl2CO9EeCch
YUMhn4NLt9/vdz5UKcQ1e8+ScdSIWWdWOEeyN+qlKRk76Lb9a+aHU87j5MSejsCS
3oGuRLZoQLLcYPlnX9VbvTEBblWVliYTx3JAA2bRp4h3KivcKWt53/NOusGvQWED
RETG7x7ByNLiDbIOVkpkh3/FGBpcZDlOKVrP0wr0MJgG7Eh/yfK3sOtIahik2gtV
9UDy8v7LypuQuXrmLeST5xGlFViUUmJAGEAntjmV4WddiP7yupNLZWUAQ23d7GZu
btgmycdiSjhkixnZUmzT2/AtPIwc7lA95mUCEQogDXurJhZZlBuxDMZbyPML7hNE
oX9VsMiE4DHzyTtBtvx4ld1Q4vmJyWH6EGC7AZoqnCAE3aqa+uRTDhXdQX8rh4C3
N0AspqZBX6d+dLtYZ/jy/Y3jW1a+hnQkboR4tUMvEfDZ8M3mSXwkA9MYVTV6uP15
dl7tDCyikoekJv3U8Ev++olLEo0jSxEZbmAAB661oaDrcfRNTEt2q47pMeTZLRGf
Rf8Br9AphxzDoJC2+Elv7VbKbQva8MiKZMpSRikEMRcYPWUf3s6EXqw/cHe7U+TE
h26EsmmazWS+c8cNEcCzF+nvOpOFwLxYPwtQd20Hzt31ZNog6OMJgU6JCa8gAYs2
t1KXeI1Pci+xpLtnG+HdfiaKAn/xofbHbk2odTYYg/zYG/FwPIuOTYOiRKxAnRoH
iU97KsXhCiRVfd9alW6abZ8D5xJHRhOq6SKCX71OJcIeLYN3KNL3bTWtIW0TMZSH
geMj4MFC5GbUcDho+bHVjrFb9ecrIpWdkopC+HHSuS5oRNHG0X+aJvIAfFbFjgJL
25NqRZSBEHl0XAecJdCE+FVb4R4611NBxWOjAv16uJ1uFUudqglZTS3FX3sh5NK+
a2hgW7MJabzmK6EvkrAlnz5cxqvlrIPLqZzuR7dZIfY3WlEV+DgZGECojPsiY8DD
r1A3suZaE6WODuVOuyV85375I6eKoQOqeyEneLWFm/8AlgNdtYNpv58LzWzqtvyn
LjScDoHqANvQdnXLvXtpQTaEZoMzM9rXCCKZAinACP2O5TkUL7JHvLFmDoAr3c/g
UefnH4QHBXlfZNGHlcCyNp6z62h/SZ3y33O5jLXOoukNqmhbMEWMN9um575Z6EVc
o6rKv9sv7U/cI5kCkIjtjUAolqcFReI2FHk1YkHPpjblkDsPwCcwwKAe6iENG6dA
fNAlTxiX8ScIE51LMp+YllKo4BN3e2K7Inxfw4Z/1MVBFkr7H6yJCAJ94pR1fEoq
xpPoTUyy1isFIqOOC/ca4066nFLEpnaOT/2cSB4e7cmw1L7SxVffRDSE35mgJl37
+Zzlp6nhazSOrMbHzYtM6WZ8TIOgomEsMtWQCvtwvMFFoheht/i1w0LdcF2EBIQj
nVLtBQvWDAysqubTsCeow47pUbOrS3XNgpuE7mbxDztNP6sDru5VzG5RNSfNaGc2
vm3SJGVUDe4ulG1r5GL7PZvlJq4I5lHlMQXTJHDTmfNBiwOxk2TH7/CVlw1TKq0l
AzfZScoH83eMscO82ZoCFYyxMNcGRubH/XoTNUlStqqct3zuS9BPvUC52qO7wNT9
x5Yp/zrBQgvk7VXEXiCs4t7WivK0A33MQvrZbK1K/bCEjoaTVJqGD9gG+gI8jgiQ
0eILDAd3MU7akfdsMqE28DOWyY5HVBsGT1dhf6LuLP2nsROWb7Hf3eLSpeg1S/12
tWl4jANHy4vADgMieSadZEGPKYJfTDOFGDWn9AyHr2u1Wm9Lh3Qs0L+s1y6qX7/V
8k7Hrm+6jpSXa0gND+ljhl+VHpO4Xq0rLayMofxwv0rP27ZftjwKxbuJq8J6Sxbx
75aS217jn7fLGA/JJR84xFgRfvNDfKuyZ/TKawropd7vQhFhYPPgXrf9IAdT1q8u
WALl7oEz43CayETkFM5v1KznzL/5IY1SkEsHt3teSeB4QR7GWTguCaG9qFKIp0gP
ZhcHHPCBpJt1iYM+ZP8F3Pil4SbmiRDVAS8FFD8N0yCK5ndagavBz7zixzL5+wWu
kjZ1oEZMZyA0peodAmsCGP5dPQgqK8jkgok2J5T+/mVvOztqG3UvHKmBK6Lyd4ok
C8haorKi8omAv5FVGeMvpSF4Pa/2MbnEc1USx4o2xuthlDBTj3QfquCA+sHi90pK
iCyrEF2LRIe56DrgMHwaVYVE+TEe9vUSwhAOe44kRpPYnXFj7ajGy2VOoZxFdZyM
PaEFOey5wDEEjQKEijMQdYxVuT/58pHAsr/IKBop9OqUpStPELSgnpWwFbvkXclh
FohJuUAH8+GTyXib2VSLzAr5K1X1hu+KH1VxQ1H0GmZ4n4R7ypCfesbMLMfejcgS
AvE47Q4RuCxPtluoNVr+oUrJVV8MnLCnccto5gQHKc6rssVWaUJLi7EFV6tSZd9c
Ez4Pkyicqi3sCevzFjnLTy5E1ZtlPFPD6+5vPlgWwly02qZ05RVFYaXFlnAP/mI9
QNpXY0u/7cP1IOGL0PsGstUmD10f99HMa1AT/XMArUmAoaYVSqlAd2k2BRk55+jR
3YKCJtD6UTrHoIDJFdKc7Go9s6HFdCVwKXopJ39G/95HUIQUf6neW3oLFyc+cBI7
pRk5RsrUvfj3eQvycatgQEnhctHQBsqmvXM+RoXTSiNqp71DShqMbd0Vjg1JIteU
oRojRTCtEm69jjckSZE71ZROj9KJsg6jgInTT3br4hLb8FECOpouisZKPjzr2pU2
8HhGGVydYm9ipMwDI7C7AhmIJXvsoBgSjb5AZ1H9lj4tZawHMsMykrXMGpUsgcaL
a5J3qLAeNyen2JC4t1X0E4RIPhEND58PKPliiVVsiy/NMUd2RiAv6ZHH6u3P0A6m
F0WH05h6y/YB1q5hlxnoCBsrOhD0jC1xQ7WU2ZQwW1kCFyK+3WQadrBuw7XyUWd8
WkGvdI49mvK0WG/W7IWOrkv8xrrVO5tIthHKX/kCGI4/uBx6GsW0Vrv3OcHeGgMv
+0qCDVsbRSnMehZI6n3oq5mPoJFH4ut5DvPTp+jzqlSKgx04ykDo2/RpQ60HF8pn
1gBX6w1Zb/R24bc1U0hdokcZeQLr1FqRRU4Aqo/DfJq7qZ6oHXHUQx25Zo0SHRRx
vxRamQ+DHkuyx/fE4SSXAGgTfIFAWeaxDdiwxqQyuhmNCDAeyHq3dgdP886l64R4
eJZ8nLiktTCwnqrkukzt0bdGJHilsDgXDVVVt+tN1Hh9fxoSKsvxk9qWkcNOJ8Ze
gWYzEEfiW7YBXuqD4IkqV/7Kb4qskQSkwrUpZMrqayHgQWLA3Nr2o8wWtXBMnUpC
IPbpLCK99VMPWjWRgLI9SqJOEekmQ7YpIst/Kvz96qc8hd3RMDM5Vt6Hr2hqY6/g
89ZqFiif3j5nY0pQHF7DUZw9dw5biifyPtCP7hJvLaZRUzwU+p/gJEezy20SLzRf
6K6x9QzPFpWBy17L7MvOqBCLGT6dq7b5+U+TuLe1cB8pYRWAY9DgeF5LVIBSDCi8
yR11qEP/CVWhNCveoJtyLQgD6varW7n6pB+8uYc9xUi8RnF9ezgtOdKmDregaR01
jiN3Jhnq6IYEaGBnBAtS7JLtM3nMRflIx2LnbvDDWVcbguWM3dYx2ShUT9aPRN8f
5dCDb9/Tyq8xDhPCl5AxkeE9o/6emQsDE3wnYGjJiFS/8pKfCWTbRrxYLdZ5lpsv
tJQFw7acC80cHiTLRNQp/jVa2pwJDpazMgzZIDJeDyvNU6BAgQen8Ur9MGXwtx49
rjTPAMWSNPPGEVhctbQ2TqbLdIPn5J+lefzzX/CASGxxDizT7T9iZWF5C58XuVQp
us+qMlyo8dAd3Ym43ZhAxfsD4S4UFx2Z5N93yBoxEUEQORhNa+exna7h4bHlRSmU
XZlPSCFe6tBZ48V1RdC75jxjWJLo+5ONDdEeAq70/2A8RGbsnINVfMgZsWA0K7FX
hFMN2ty0yPhBqw4MVNDtCCT3maFxl0XWzep3KBhDy7FfljHQJ5RBKwN8OylGiplq
nByxPqrPsPJvs8Z7eQqRZau93dTm0VZx5IcnhUf05oLACUkNm6VVkQtvgrZxalW7
+6hp48JybofwzelqFeK6xCyqgycFrfU80APYo90KJG75Vqhlc4nI0TALKCq/jJyW
E30hV+4/gGzVWO0tA01+/VRwZGE8iCD2xYvV9VuSgOevSZqtYiSQE8YXqfHNp5YA
ztpHdFal1zVdgydLDCAA9wwU0P8X+T4uQqFFk9WnuYyD4O6CC71zdp4aAxANrw9i
EbvIIl2QmipA/yJzL6LeH7oym0WWIuIN/ivg9XMi1+Re0g3oEiBWnT7iRWaj+WLv
Y5o7L5uWnJwpr2xMBs3gK9kbicukXjJ/gtlfa6WjPwHtbetA/UeclUPW5EvTqREF
Cf7Hd/HD1iHqfEMArWG/fCkxcpRyglO54N0YxpA+QM4lUE5RhNZ+vT5AROb1rDX7
Yta4MmnLLgefWbZgxGJX1L/HeLrGd2jm/2SCRX9d6DCarV8sPa9v9MCOiKYo3Q/u
L9fsMvlRZm6eTBCtJbECaR49esycMNx+pfwvStndlOyhMoy6sB5+GtNKoAchuh7j
kYzVvD+20VyclBw8JicqTZ8ICTJj4U6OLD8k4SGiMdbVvEyYtCCuOGrk+D6w4iGP
QNpKgDSIAPFap5CeP5P/zyr6RozE3+JVIpAcxOSCjIWEH1JkuFSkgoscsTO/7krJ
qd95xTjz4aR4pTLUa8MAY7sUFCAxUmOPgWi+aKl7qg87pc20ikS1RuvlQ7lRtSt7
vtGNCO4aTa9vLP/1ji+bBnQfkrBUc8viXVHCzbYygJLgcdKPF7JFcczdrt+2fqP8
VIMM6rjsj3RtZkE0GT9QFCb0U7xOVQcHa2l9SyQUEqzwRnCZKmuK/6ZyUWSOKZBQ
e9uQKk0ofmRsClNWNcFJbOJJ4Smc3yloPvZ5ij2Hb6oyJBShj1xBrV6fUgdWzkeA
iQeRHCYZh6FqHDRCqcSsOSy6HnTK8z5lODz6gkgWpWCNrP2K/aUODeKOyGtnGMgv
IEi7jdyPGLsjcviln2tJHefszVqcsnjOXnZu9DC4i11w5L4GJJxVy0Pe/4hfEz3k
mMsBZxrZtuBpuRS23DoAemgCDZq8LB0SvB5Ckn0ZfjNQFqcPfzPTWz+KOKW/eK67
ej1UgD4gEc1XU03ezlrVBJyfcClaat//gx/5/YemN7nxrLYByuf1x5ERd3ISKVu5
hSWQ41PMFD+X/IwzKySGlAo7UA1rs2fd52qsTVVXpSVHnb4AfK97xS6UGqsmnc+f
fZGySf6A+HkeP090Qt7wz+TzjoyW2ILuEmmjsguNcRO7/VbbhkbJJBRtQ6axJ+Yk
zPEhyJCrdDh/+1qPw4rLK24tbgK/VbBapG438irWbVHkOyV6+eWraDDB+fUqhbIb
mkOqiPKTc7qDB1Yp+cXS15dlrh5tGoXYAh8iDZ0+R+KqNklBme4/JoDKsaSX9JSj
FmPyNoLF0LFcQVrOZpgBSH3QpOiFizsdZ7b9UlLcxTVLTsGbd/dq0PDP1olQKNSy
EUB5n/hAJ/M7bZBXX/idMFzFlcwIgUsJHWneV6SG/ocvqf34/1XwnDq5eU7pc9lm
rt+S4zz16L14OuCO6p3obQznkg0MMyaGygHUbiQHjhE7QOnjg1BaFUDcRogXnCoI
5QIcCyaOteA7VGtXdV6vxEGTvlawpIhcCVoF3KZdgXgBBm8JmVCE0PEzsxPntqzg
2bKd6b+qnD+Owff+1HKGbV/HH+cXBeg/TqZZMykYL+oaboPJakdJZdZuCU8/e79m
pstO5da7+RX1jQYvyPJr2ddwDT46eacoXzB1oisOyh36t5say1fKduNmffy6loTl
O3VGyF76krDQnvA0ADAtQzzy8P0g1HSzQgcZDQAiKl76y8mCifXV2BUqXLp8WFKI
Y+sYVd0qqto1ivsl347EqarDhHy0utJEm1yZok2uDAfyf1a8m4xTUMxtRHicMh8H
pDdIcchfAR0nF/wgxZHjsZNS+/2NtmacJoBO60KJZ6sc6Dkf6ytRJJ+t/tUNp6nM
F6LnAWKVFWJ6gkbi/XIYh+RF0K6lb7yADp/wi+nqMetePfc9qJ1BTpBoJEcDqqKn
q+oYxG3tCZZmyXodeUFaKoQ/2dBeFf4XlPQ+KpFYtiO//9lCnM5bD1jbDmiaPWJo
FRpxd9MNOAOuD0nQ1hEYCujfuk/UgeaB/l8NAPqmqI1+HnUY2EMxON/Wezuwf3lM
yrdxnhw5YP6It4UrwjvBDqoCLQnYapuV9ItgWGbJzjlsAvLjdAuy4J/7ytyxzH9v
uwFcuRttW1l2q4R/hz4TVvI+ivxSmfMa+Zrt+pfbN1Q+RX2XbtMyQTV+jomE5Vpb
DZTWlTp9ds8A61qLCAsRyvwE//2oEjCcaZVS7RHTswtNPAVzi6AahUmNKIXScuCZ
XTtz309w2bTL1/TqZNRVgyTC0+RFF7Mka4/+DZB0u8pf39vLd1PPPvLZ9qbOARws
Jt+q2Qi/A+uBMi8NukcVvgZMzB4u7xkJQEjgb8oOAWdBeuiWd3DIz2PtQCmT1Pga
eseKsgi1yeCKti9Q55zW+aW8dNwycf1/c++4PisiW9a8CnO3xVY3rpDdJlQ91UbZ
o2UNXuLdCaQ38yAC8t1erXXKzNrur+1qUk7t4SIIoQrDn9YQs11XZVcTTcAU3Eqy
avKV499BcdSnOubDNkYjxZNw6HLWufFpYSZZULwfut9r5EEL3Oq+69BEPyFJD7j1
11y9Vyl8/KB7FTzbLXOUFivdI5pcU4NKKKMzd2IbKAbg0diEmv9n2InQohtkZE5O
WmJBfQUi9y4AD7IH8zlMunu4ZLX/ylZ1W52pM1FKjYetjexxOUmsgpnj0eDA3GWV
aHy9BMo5XDtMX7LgX3dtymYv/5mtjjDLrPA9dMQ2GexeetVVYUQr40z9Yy2VXNlm
wV+fYO6mfL0i1pD5cwGG8Q2Y1+1AZqSb/iNUZr6e5HVM5T8I/7fHn7u244TWbslw
LKP0mgU+IF2lepx8vQZEqswLl80+c46T7CkEXTxi7i6P3+2Daqn3tKKp3GRAuY0M
CZ9GMFh81xhZpbk4uKpoB7tVEqpdtgtk+jLUI2pKUQltCsR4Gy6Q/eQRlUswnim8
6cYuErJKg2JFH8hI3hw200gBQ0BFRMLfDzwmKQG4/p/iiEAuLXs/baEYSizcEDuM
WACDyMtnZFCMs1yAQ+mfFEFUUCaRVbW5STmHQSq5tNumvdCA9vz+Vr3M/PWQQFM8
E69I4JVhrEbZ6zpYWt8R6DevNBWOgjwue/Zt+dATm8+YqoxmuYg3N305R8ACcuAg
VUh3HpJEUrE/FTNGWDah6P6mOt1xCcfPd5efwacp9Bq3rflY82/XSzpsDlveRuKW
+vO/a63itjVyLuwwpN7H9iSXFBy3RWMU31FSt7NRPer2oiFncmCPOAM5jQE0dHmf
MuTRGQWU//S49XeI3IcH3q5zojuydwHOLbcPrD0R3D4wVv/rKGeDUGWzSTK7DdBj
lj84UQMx32sESxJzzZ4g/IYv2AVNFKBY113FW5WBj5Rx5o664MUx/jNEeYg6Qoel
lZuK6iep3BWbpCGMfWGJQLbiy6H6imnjghAt/pkCUoRULVPsDreDy9tW3iYFYofx
HxRQRhNkBvc32njAk6uXr4j28VV3BqHKAuL+qOjz5mRJBflKKfprso+Khwh1JsBo
OKP4bLwI8npEWAf27ZQPNUmWA+OU4bFMFAqfm57uETYmE37vmkMELObKMa6uZpxz
nLhXpD672RQu7HNR4BMWMra8N1iUIEMv0j42kii/Xu/vh68FPvH9Yxvy3cSJ9gf6
qqNxMegKHb6oj0wDqIGZc25vuqu8lZv9f0WlD5HpdgavVK1tLL0IEvMKB7cli+ou
V0iZGGsR1YGDzeqi+fjVb4lOQzkzpPhRbeV5sTZaOunTUpNPx8RYCsnpo/D+Wjtv
8OMYpFPPc85mhcSgBS1zKTN2FvASgkCpPE+WPlA185fxZs1GPKq/Jle5sSfUd80X
qixKa59/OaclIuNiuyrmTm9MHbL8X+eW+Nx5whXHSNQ0Hd64hJL4tQvFz00XFcYf
RMaeo3CTXSm0i6yKrEUqWbdSrMmdaDhFi8EE6RkflE8JHluD1GR+7gvU6gPQD42j
566sLDetY8kL5B9lRzzIut5ONbTqwc1oDk+Lo7oatCY2I1e/zOan6IqZrlzgTEXS
u/2PSFBxE9S8AIhnr1+g9iW/bU5rKrxdUGkS9h4LkWgc/yR1qXzBfs2HEQjlC3gu
FaFDkwW+hf1Prj06Ar/J4Q3jZ+ADqZETn8/SKIZrtL93Q8X92h0/TlZgKhbs4hdg
A+rdx/ddpdbt0aE7G8SheYqPsVX7Q8YkXsBhoKq1i2trM+GEhwLLynN/Ep08b3cu
+X1YZkXtP378wKEeVq1ughANCR5Zn9/33pSlZgbLKQ4SZ//aSuRD41HYtgL8yE11
JOGYyBjnfNVeeDOzEqN406nMYBSS2swEJXaq5LsprZ/0BrWXzCKQv5FeCsR/+3Ws
6E1l6bMeNxMcERR6J9We3e4l+ahrZ8LtCF826VHp/JmHmGTePsgR6zy+Ir3RE1l3
HJSMud2Zcs1uJygVrgl7UX9UfzfU/8EkE8D4Ug8XZQ1CN3sOaZ4XVINfo5DG+daL
MGCG3InQ4nVaUCQWa4A/gwTWYKgtxbYVtlrlo2W8xRR+Hjzd3rYSYFkKq4snEBnj
ymBnY3jelRA5TaNNSOZ/ZR5GWlHgpvbwEngHnuG0BMiXSQ0XnXtS0kIi8XZi/HmU
khvk/3y5KvTW17VgmjyojYONtSpeyuj0tX0uN91ASJqRc7Qhm/dsqeHC68PL6fGw
tXWgImAaK9rLSsCXOeHgc+UhxrZGVOkCngbQ0thQdS+QEplUCL/CmahxPFiMhyWB
4gfRAzJtZAGv0xPgUGyo14+E5uvIoLWQaWJ6r6F3TjbIgUfOKWhNq2Q9SrAU4XCe
WXY5ph3E/umRIWeRATUk9slf4ZcUKIFeZzWB99mrrTNfYL6hdkuMuLLXwI3sIbQE
/a0RXpLKeZK9iMvUgUHEYm75hKlOWhaaRo0LBe/ybhig9RUkKTxKkRxIU088vpfC
KeMbf0p1Rb6GTzEwmfoWw3+YO5WBwFFfqq2u4EXFaCmjO08/PXSLegb9KrxfqCQD
geBGbv9xkMMsOEzlelMt3WFqcsYv8pX9JMBQtMUr7yGfEcCXA1TDTFDdXX1M7q/p
BBFRJ2WbOLoxlY2Fb4GwkA1iEO1/RKpcp7bLMfVkks+quTcQ+u1kXPHsP+1cO7HX
ttHPOvtn0rzk4TyNNoW6JTbEFJMAuKl4t91as+riCval9EQpass3nnxRlOpxupNv
onGZrZ6G8XlF18g5VeBu97cC3+Tra8qVyHSxCrs1eepysHAqJldnc1+OqSAKR2je
VGHbI3unjNHjf96oWR7Az9XELInTpc7DqWPU5b3QgjXt+Wqks7SeyXusN4TOwNC2
yGW4hRWwZjU+f0b3P+8D1U7S/LEmT5hkU5aY2LugZqC4kJiclS/gUEnfEwPA0XZV
Ej3LSeqoE6WR//aOURVZVAdXs9EcZVuLtFJSRZXHSVzZ7oMHeH/UHo/K0hCQLARY
x216qq3MkaHTH1J7UDZdlc40fGBcuUZIhtc3KEF2l2PXPjiz841YQ2tHEp5VR1jg
6NdmqGt1I0xTkNBEAR9ZhSEetcm6VaKueBibXTzqieju/E5FAwaLed+51+a601ek
KSzDCpwmWrQ4weCBvgcZq1R8tzOqH4Vy/i60383y/pq0ZSiiU9rYHrXqMLofVIEQ
mB7mYruO6xQ7Fp+kkkIIM2csXAHgdmnwDNrCjyTA8dAm4sbWLVTr0m4vQXZVkVfG
62pHgUqgD6s/gHSgL6l/eVSQaIf5l/k7QtKpHqkdIR6R7uobNqMRT/SUw9KtItXF
LRRLy+ZWF0589zQbjGFUvNC1gLcRgy33fIQK2QcX0VzE9nqAUNGU4padDGhS0kco
mQcC8RudxnP7Q2YltuOfpTxXz7JA5RYiQxNSNxtExOS6x50B5ETD5BYGBb5Q6GL2
KhRdIpMwiI+zFL9rRIK7WsJxmhqtrpNE2vTsOdZRZYg7lUNwJdQJNYr5+IWAI7m4
1c/dUNRzMbyIRH1kkY/QcHlbV/K2ixhSaFVHZkCw+ZedkBBKYl0CEer6oNVohMM8
iir+/PNKeyluZTgHb2TgLx1Q6RfBZ/ivmSUFIUMw5SUf9620gsFGyyqQeuqx+2fl
in3jXHTCEcy2fGi1FR2fpaddP2rih/xT5a37t7N21kcJZR8ExIDh4bGdgMCnmU8T
9xf0x+TtBbucIFOHspfkJc3bmV5O0bXJrPqwc4sr+yVLFlXDzgRuPeYRwx8b5hZ9
o6XQm4EN6+63LXCmj269VhAyszhujJBwnGSQ0zCKetwqkVwvs9beMeOXBwclwsWn
lOnNDSJMtdB4ckUgSP6dQDN/sPn0OnuK50SrQQwZq38m9+U0yrEpk9kibyUKGVlR
rOQrNPsZ6YGBPQ1Evy8y8n6eyBqOUxDm+ysEn6gtF4cY8g2lLyz7EuNPT+IgShWB
GB344whR0o1Wnc+vzYf7p3GfTrRR0z3GG3VSpdMcgZziQys0qINzX5Y0TBA+kPbp
dH/9jIe177Tzl2ThRRNs+eXFrCtg4ODpv0gG3gFwLkn/GoTJ1pQBjN5thLW1AE2F
eKIq02XsTzYeL/P9ji2QA+gzEo0EkEQ+JHtEY91u+x4XmPo6qeLZQ3FpaUx0l8uw
ympkai943F+mfun3AIUjaufQuZt6xe1a3jbV53BjkkDyFRZVpEGr2Rcl1pAOzCgr
+/xTwMDtLS2cpKLUZ75D+7skApCCm0GHAl/oNmt+GQimR1azerJaQV8Zr1pTiITf
5gF54t4iW1+nVBPp5bXWuimJJLALUiIYKsmDgRaktstfXsvFaifhAB6gjVm/lFNI
ywSdLq/mBvnG/4gT7nnvhjq/MaGTReT3iqbkR1GnJlJNwQOhQs37Osd4pJS71ydQ
GBXrmVXQo2OOjjFmBapzrC1mgi8mveeR9FyHN08FcTElgNQY6XswC412G66umHp+
IjK1vvqkpCXF1pK1q7r5RZgYRsyjhfmStKcdrcWOG0LqhXPsEcbSUH+qs9ZHCnxt
+3Ws0bdE5bm2p3hf/H3l1ExkOC+e3ShxyamATRuZReszxvXqUOjsDGUyBSNRkop6
e2ll7xNpyXIV8LUF8P5rOiIcR4T7tG4zMgX2/22Oi7vO00vapuyN5FnKjzTs6Fly
hAEkXOXpC7JZPVdWs8A2uhRoE5qmY1ZI1kH/YjL7XMtGvwgo57udPIQvtVzhd/x8
kZFM8SMyCe5kraUgtp0zGd1xODhbFxGEpQQOqXC48yOXpaydUkN9jYpw449ysz3n
wtJcVDuzoEZYRoTOL4LJod1rzQxT+VtbpMz0QCARBGIAshUJh8VdPgiizG7qJJuM
HxJFaovIQtk8vvUBa61Vz2FXP652343dtgY58ezzA37uZ1rlO28FujLEkydDsE8X
qXm8i+s8+my3H1+9gvJcdKd3H3PgUq23NzOXXY1mvN9nflhfnRbTQl3BZg1mHNGt
U9RGgT3ZTeOccqGloBmhoUA36eGUwi6fWhdXLobj5U/00dRkC4SpgHlC644E9MkK
rfzM4RiXDOB+b0cC5kdahcCrFitNvdKu3mgG9Kfkp37v4mTLUIB1XYjActiwWEi7
M5bkSYWA1pTCBg4akeyDDkAOu9Z7tPQ7AyE9RVyKIoeXa+HIBA+NMMjP0FZueaPk
dkcxn0BwhDcvYcBSJVi3cHkEYfW8GUEMrFDbmBeEv3+LFUAfyF112VhLIHJlNd5Y
T65YP/oi028HbYdkhnafS2FZbuekfSYjOGD2AYTt6Vw2TRDsHAk3evq/JztuzOM+
2GNIPiish2lgqC10/dgJql4lyBL+vNer6cyX7iAJPGKo1AfKyXtXd/Lf533xsq6w
tHyGE9L/i4qdMGwaZt75AhIMjYm26arBXuRlu2g/gicYdzBlO32EJazubqCSELpP
MLqWHtlqC9GCoxY8qvrBcjIImtg6iHnF5Fbhjlud6wauxnyxTPzG8ZnIfaLuGMx4
KItMbPLCNclXSpkZM7m1zVf2VBE4m9mBRfJWarZFHpePkKf3nqxsNqBqGYuaZfUw
GG7pfEuFo2LiWUxvDv8QMaGEI78SUoqjxdXA6Jd954blWT6QIc99H6Zyeg4KonYK
eP6mznjwTy+COiThW2POhgaEMrjAB3v+8iti1cqI1hgBtViZulMAqM3KVOh6FPK9
7EQQbrguoDx+2Mhx/Yqp28R5Y9RB/nUYE1xnff+MfIsLUqvFYrr2LS4FIbk8+yKw
JLoBDqW/QRIjOhwGjGXFdc7RsWSGXemGpX3G2dTv6AxWRolNDi/UzDs923xftBQt
0H3F12oFK8xu3WQCt9ADnt7cn3PV2weiJp3S2PocJwkEjDcyZbQ37wakz1vJs79o
umWoyLvrT5vufcO6M2OKSPTpW9jExx39am/sKusF+OLj5/DeJ4k/jzPyzOghvzAw
lu2/2XuVrE9rQGK2t/80KuHSZH6gHfRfXAB0AdWj8MDsVXl1EPifjxGUWGRuhRQW
+oqb9/z4IfxN9/cQy7ElIOMY//v+Lv/6eKiFII/mDKf+Nk5y3eg9Sw5K7UNGKR3b
WR3VqufgHvBZUksY0CLsw6C8vKfJ4PO9Eybxhhy0vePmBbrk3rig9figvJ+Nqmbn
KCf/+88rncnLeeufMT9PG4mxWpF7jggGTG7GkMhCLLVcM7yv6u3Bhw0jAKiN3Waq
xJA0KMT/WaQzND6Edsi2sYuE7V//mrpRomShNU93bsF+2Cgw38jhcmQH2ApTVIs5
PO6dUfwDOP5obteRcwDvrNLgblh8An/TgfmBux0rt23vl1szpZiASXPrhMAG9JM4
fBvgXnFlA30aHEHkLRM6T66vHSx/v/A0erQPPFAhqvZIuBx/4waRJLYzWDk6BP60
Rp1jcezhsoAiKQbZMKrUN8Co8XBqFc7oGHMGSnDOB66iSWMLwN6fkzaVyZn5RL3X
bs3Ksn7Su+or/+VXKIX6mOCOqUE8WdAzxDmhNgOek9Ps1aPGIpJPSs9w15P2JodO
oRN+Upjq5ysOAvlKCGM7qFuWl/9hC0X3pgG1j7FR4bHK53Hvdtc1laja6a1amTuF
pkNTDWjitXjga6ihx5Z6iKWWW5/T2SpVARJsFicma/peesb+bHpcZefzhGfdctlH
vhIkDi/oFPA02AhqiDeAD6TkkkGbg6L9QeVu+dbMfpYua2qSbxgOiYWYQzgQgtCh
syuppEXzu9c0ex6G/2TTL8A5qEj8+3hYCjHJIy/p8bn3T2ZXwze2eNaW+1YbuwBG
kzo+s3Vb3or6S7nyqSMeSyV+SEraakXFLUn61OlV6nH/dl+ZtctypD/eyST9esZ/
4i9C7gbL0CrDzVJO1Qh732CN9189VH/6F8Qw+R4lfsnx4vy0YeF9Os5ERThLNWEx
YDXjq5nCFLsbEyc0RMuku5TRm0i6hZ60EktQprj3iHVb//Lxmbh5lRYX8208ydaf
/9HRyT8hb9yidthlApMUbO+lluq0q/xzhbxr3LLzLBmrQXDL+fgTvkAS72K6C7ST
E+R8Ar54nfNEu5Bv/GOLf5arptSw3PolwRxkd9DcmOIFG0qowvLnot0DfVLjryEC
tHfcauurQ7f/JCR7w5zoCR+1cFBuVYMj3D1lJt1zLaO2TCuVOBbSIl92RtbVdt//
KWyZ9yK9SNEuJBsSY7H0T1p8ekLyYw2mjqrRFzVr/nSnV8yNsJYUpCWe1qS3L7yU
2RKnMYN77movmiUZET5Tml0TzIGQcqqSeEz5OABujdVbQ0XNVvJKzDYG7g9gqktr
inB/kkVh3MWRFeGBmw/Nn/9lyRCHcmt//ORkkZMzUjD7U0mP9dTxSHCmW9JjXPpn
JJ7mV+jXLaGPmN2r/YhgH+n4TXudlsxy2lFLg85TqOYl9FrpqvIuRreRfUslD4E/
6p0aqHNBXkVgMTi3VOZMFhA8P/FLTJxhDA8XYuE+AXIS/OihpYr93hmhISb2WP4q
SR2H94mMWFvgJ+ACpCNsXahNLtoyeNA6oZskBRTmKROV9jeS2Jv3wEDx6a8N3nd2
tANtAKPj0GkH3sliaMtgMOwInEhHkQhRxIxHKiIOehnLGAbMJNS7VMhidaOPDAR2
SJvUBxhKkMsLIl8p2dBsF9/x9GxqNAwKWPXscfNKviPdvbPbw2vdGHY2YEHTCU4a
CuvnFG53JncYdgtv0tO+Q5uwZa0aXT4Qh/htWSuL18bGMxTupqUdOK4C0kU6iI4Y
RtrD74xJMP/31dMU9C2+gol+hKBb0zBeaPEzBV2uwjlDPBiWL2pOMokGvaNMg0vC
jzWJZS7d8lIDKaOIlADIzSTfQDCJoQ4c4rmJ5qPZps1/6tGA2HWKCtlNB9ClYnoa
deFme4MC29BQQtmhPiSqVAQ67BMr4kwdGau8Vi8NX+I7qY+oQzRZjqldtGLe4z/o
ENAGyjBmtlJm0xlJc3IGYktdlSSMkVuqXW5i+VcIsg0lyJwG0s6lrbxtLSNdi+lL
r/gIh3kvjgK4GZrjGEqlS8f/qDfNQU1sttpuk0u8KeBzmss1lTPWQyDaxcbQaD8B
t9bOik6zilrjv4nG29F1RXeXWZfAKD1pjL0mgLFFzfcetY5L+q28aLjWGH1It6oQ
0lIUEcKZsRKbgZW168D2X8Gjb0mnNnZJgV0FoE6bBcA+NUH1YU/ayVrL6dwYDugp
QrcN4+afTj+HqKPF+yPGxxVljGrLTn0niPtEsYpsy2SO1EbRBTPipczmP7i+YG5M
SHPxG+OFue7qPFKotSXV6vgSdMk4CZjNqBeCRezUGF+vVsLBW0NhUjwujcaQzj+D

//pragma protect end_data_block
//pragma protect digest_block
7hsRD+IOdtdxUkigiVbfREcXeeY=
//pragma protect end_digest_block
//pragma protect end_protected
