// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HOI;")&M+KQEZ95!-3T37 _XDW'9P7?8V/07U X\K05'^I&S^\+5OP0  
H^@J_Z#<.:/DN$HXY;2>RR/N"<A >>EW2O0K%X]Z%#.?K<3$Q@! -@@  
HX/=NH#E'+JF<>N''4_U\9[ZGE)F!%9+\;+A$V2%Q>G'3%-((:-+Z@P  
H/NHZQM:"/K>7.R&W+D6JLY!XJ.MDVO[>U,55F%Z1Z0^LVPX7M,1[L@  
HI?2ZS+[5MW@:\T%&Y2P],M]455MO#\*D=AB&'58".\%N<<M(L,8B20  
`pragma protect encoding=(enctype="uuencode",bytes=13664       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@$ZU&4,1S]-L/MI%1*00=5(\1@"F$3L#*>>U/;*OJ)GP 
@P[)[6(7LTON<H$M=!Y_J+C @LK_3Z8.K<-N ,D+I"^8 
@T\@5AP&)@(XJXAH!>8FWSXNQ)J8&*]!Y7H8\*[6$_9H 
@=G1FB&._2.-1N0MY0&C-8;HQG[;L,$B.\.D'7N65<AL 
@E35K:\VJA]ZI6B<_31NN7Y#215K:"T1]'B)U\C?O@L8 
@A;X]46L%E"Z5-D=!!RI3?Z&0G8;[XG?@]B5JI@U] 9X 
@@_XN"?T>KN+I,1T!9?_- []#PRIW6(A H*4GS;U4@<0 
@31E/T0&L(/)Q[@=!^>0<#1R2;W# $.7TYU\3'*37?@, 
@Z&DB5Y@O+&M!(HT"V4[8FR-+1A9@>%'@P]S>Q4M*$W4 
@+P?,8=*G:<-W 5+ZP&LA]?K2,6VOH0"-F5,42V@)="T 
@QX(- ?@)DJ<&)9SJ#<SMUL-9U6_L9#*"F[7H_/-M=8L 
@^!B240V+'->"))S$+>RJ1Y>"F-R\_08FJQ-LC#NCV)< 
@JY[O$$PPJ9Q>93'^@5@_VZDO;-0:3U<R7(3<9E)!5X$ 
@NS%KFMY\<4=$/AN@4O8@X3=TG5^EC#JZY5692W]#IE0 
@>UC4,U2!\ -,[/ANN;-%Q)2&)]U818L-&I*JQ@<"JUP 
@8HKWA2(5>'J)UELA+>-"7W2M71DUL\$K1."2K4X])SH 
@9RTHD"56E6(!G^[27!![O97-4Z"S>TQ;)/,33(!LE=X 
@0 =@2<>?8P T#OT4YXK=/-,:&KVYY/#[T>"FRVX\.%, 
@10-M9ZJ+,US^$/33FEN#C7P>C."TG2. :;Z"WH;W584 
@ 2#I!FGC:05Z/PU-MCM<-%8)#Y7J24;9O X#.T#C1IT 
@'-@"[CDR775N3L5%H*2NJ0HGGX*G/VC]>A0[>H^Q.<  
@#EX:S5%/&T'BIGG,&O=S3>1>(G]X4^U _$?;MCYLPVT 
@$G$5"<7DM?RL?T6,2(K4/^F>Y8B]9"-['O^DB5TI*IX 
@F5R&=G[N)H7LSNUL313;#O6HBW\A-;EE_EK?V.;0/G0 
@0(H(>&0 8O&"AV>Z]14>+/M(XG?[/'M4TH^7%F<1!Z@ 
@QF+,B6*K/:46,-;$>?19@D"LP!#07@AP,BF-CRVY"G8 
@L3OK%L?I%DX*V@[N*!LXNS5$2UZO!1@JD7P_4K\CSZ, 
@C$&\8@JYSR3^?/5Q.H* T)R 3[5.2'6/=_.-!#7I&:\ 
@=2VW*K_& Z<IL,1751Y785V(FL6);+'Y%*E9KTZVW5( 
@HV_W4K?=>:=ZZL<I\00B@QO*4V[N<&<-YYG9MS@.0$, 
@=E N0/X'>6%X_M<:5!!XP89,[$Y-VP0&,WSKRL+ C^( 
@K$?&"LZ-VQ]^)C<"\D-'<I;.7=Y3\K+F53F#''UB*1, 
@52^4=P69 -C*)XI=,/=*,9>;R+7O>WQL1JG[-&U__O4 
@Y=Q/$H^:J(W$,J_=SZ0'W)%A2MU@/Y7*PLH!GZ=]<LP 
@T#ZZ5>0 ]>%/QNB2=IQ+5>OR$C.KJ#&GYPF.WMW023D 
@OAXPF;] _8H64ZW'YV-6S: ;-4U+]UWG_T7;HL$J>4( 
@!,V$JX?5R0]"37JFI/M*UAD-$MW:4Z,C+F!7Y K*'U  
@;54A.L>-$A.LSZ610P_+A,W]*_8T?@P9#@I_Z'OI5.8 
@.0?\9_#? 9)9'+HTNG>DW/6W+:Z?%G:)X=X8O'GU%F, 
@)HF3FO>3+UP]A]'\04 MM!WJ.D/16/P8^\A.0Q^JU/< 
@F/HW:!!QF;%DQ)VD!"W9>!(E)O92V>8[R<PDU])PZU\ 
@\O;\-6,#&_/D;LU=VG&NYXF! BD,I3]=Y=Q&88AG!9, 
@Y,0<$,+VR9XJ=1R4,)><?I]7LQ0JAGHT.V3@*5$4(%D 
@9+7KP (!RH<#"=N.SQR3F$-P?Y&7 *WYW<<TDS7/%2H 
@F;KZ5CZ$SIN<R.@G05&&9!=1 ZH'QT5].)V^C^!MA[H 
@DZ192Z8?<L4FN!>76)&R+!'-PV)MNT&%#,:J92V?_!\ 
@TCY 4J Y[<N&=2."^<'DXM&/C?J:3<-CJ%@VW86-#[, 
@Z+B_YGV>UL45ZD@2:'<%*&GF[H0XNDW<@$NV-M]2LNT 
@]5K&4\RA92A/J95R"47"S \J34D6P+%&J0PU!W?QQ"( 
@_60N^;CKY4&ZM[?61S<;A8TUM+I.> #94EN9NFBFW^T 
@*H)I+%Y'_H.S-Z%#WAX[V^LJQ*8T%$43'H0"B:T)1X8 
@V /UH&84@T?<UZ"^K.L^:ZLYOIZY<]!V>F?VLMNCNVT 
@ZSM316J)CWKU:L(ZTC2)T"$<_!"9.#+0D?SA;NG'M%8 
@0;P!7BVZR+_ ZBVUS2?R5*O:KESC^;?'[O9:NGYP+\< 
@?1+D)P>UQY*KYZY59$6?W2PAH!GE>+43AG38=:78B0$ 
@5^!%!_D=/6XWC-#%_!8S]"DMK#!._XT;3<EI,C%XO<T 
@*T7DX</Z;%MD'LO_'*BV=(S@]7;"> $_FEF%LU>>+ L 
@'V2P2(S)T#$L1^V.D<FPH0#;+4:#_2M+$KR)./ 'A5P 
@PM?ZG5QG4B3U"0"T/Z;1PC&J28 ;IK&"[TOV%?5^^F, 
@\VFVQWO22^R'(LB%J'GN5,UM(&=_"QX%47A\/R\HR:< 
@"SQ?#8_HHVCA=9SX/J4"IA65-@]J0OWBY?ZP3W4XC,L 
@BENJ/ -8)6);26:7LG2^[/8/3BA)JT>0\]W"B%>XE"X 
@I;1##3<:<4M2#Y1 G>-FC47_TO:),D^U(>/"HQ^B__, 
@*B,,BH%W]!R-5QI?)EG8849M6"4WBMAR "4FEW6HIZL 
@?6'NC*0IK/D0S/K%_0=1H")07,5_2Y<W?P]^W\Q,V1H 
@5H_OX^R+_58"+Z#5C*#U*#XS\1A/&M'A+CG$'Y---[@ 
@=!U;>E)NI/K 2C,^O4A/8!-EWXOYK9,S4,TVIFJ^ HX 
@)>^HOBH3NV=;RC*ZX; )MBXAE\$YV<'3D"E P/4@<HL 
@E:QZ^[;W2N]5Z>W@ 8PNE6B$J !IX7>(R#$%6 <@_4( 
@1W<YB8].K4BH\A^H6AE"H';&4K$.N4JE+VOM>-S3;40 
@;B04P'.WN&[K@^5YB<,G/+\9;!H8*.,*>Z$'I48F\F$ 
@803O>A]MCB6R% W73Q1=%ZU)8@<I$2 1CI>Q8J3]))\ 
@QQZF6FKJZD$5+(-^<Q57-N.'.[09A_1T%I"[O@+O'JD 
@$_4.SA-KM21Y>3R3;3$=:3B[#KK<JW<4115T4.LL4&T 
@9I84 <(6Y>/0P]1O,G_#;X+513B'F>N?^,M4B%9\B;( 
@X3GA2ZLH^?5^,R'8%)\MNL+M\G&?P7]H4HX S,,GYG0 
@1S[6B:"U2.=<?\^&?Y%<077#(QKM(_0)WNJ^UO#3?H< 
@T3RQKT<3'"641>T4LI97*XD$M%7#M,@Y)-IGL9RB/L@ 
@>3N[1> 7;]>36>=;@E,(?@_=!4K1.J@-K/3=]56'5P\ 
@)(%IBX>[AS3\&7Z38I%;?*)VHJGQE\4S:ZAJ*!D0J)8 
@+4(FV^+E_-[,$>S4=+E%8T0!NVME\C3H A4Z1/M@"74 
@#'X,W+MU<7^,F7:&$QI>W,#Y%3MPB8WL7)*@<I>H@8( 
@5(=HRK9R]2%'Q'N<%&(]T@T$!DRT?W(M.+-;(3H$_Z8 
@_-=A><;U5QS'.X9$ *CYV8D:<PT9/PO;67%5OL:^BAX 
@'JSHJIR..GB]HD>I'@2\D^__4;:3@\14$0R4 !L@>MD 
@M/SZ#N8GO2DJ\/_"BSA^0PR?M9I/#-9DMA*>BK.#QPH 
@8(,E7,L=.L^ BLIAIM;N]$);GB#+2P-N\W=6L679QI  
@LT-]TW5+1OF\4$!*<"UR8:N7H6E$\50]-]6#B0F=%_D 
@1^#;$URV!K.FWD'TPC5H[S&H'/RGC1D: 4& W6(==WP 
@<5G_-L[9<[.EI'3QMJDO:#,@?[3AZOL',DQ$>YFMK<T 
@PVX8-V2E *=JOF:..MLHQKM8.Y^'+4.YGOJE0CY0P$T 
@2<%AW>!+N@FM:>IA?S5H'1,XOVKS<Z;Y+5;ZW2)PY$X 
@)+0[Q0\=.6";UQ8RN@NR0D1(O/7_1L*.7!$/FC9J;%, 
@;$I+_-,^"4L(82V6C+:1U2:](?$7Y/;-NFOA @TCTAT 
@#,.I"^=[ILS6D/ ^Z*D?76KR7"5:'R]"P*WHK5^A"O@ 
@VQF@4WA>00DB,O=*EN<S"\3_'][ P4J@];MB$C*#YMT 
@'_#W-;1 *\AG,JM[M[]%SM5+2,(%:"=M77W6J7O<>3< 
@GL"(Z3*_9\60VNN7J:="%Q'2VB,D$/R!:_.-MYHI![L 
@4CSR(0Q[B?:TK7D'A(>;[0*PN]H.5&(DW^H5]D7&"F, 
@.TU-HG;L'-/__0V\WW[]ZBE.B/%_,3)FG=- 46[HO*< 
@$69 <QG@Y=2I>%GKV'47U0#Z70MZS*U9KN#71QU9D,P 
@F*.[./1.XIPU2?5JJ#$K$Q!)4T"?.9&W/A6D?B%C&&4 
@ 3G!N=W7MZ:2#WG?%J,MC@@N@:5X1$R]4)6Y[H-J<RL 
@4-Y #$(J<@!\ZCZ-;D&)FS SL*D=6?G<X\/ "9@B/T, 
@F.A7F<6  )6CIW07=Z"-\33?5I57.=G3<"4#%SCKQC, 
@@M(N9 *4P"% U-<SK\RO/8M<65J(9)>&30L<'_A&..  
@A /VRT\XIC&<<;/@+X*;>7O^Z^9\?HB*5'WQ)#P8"X( 
@FF,RU5:*<424O_Y $NESHGI2*5^F6^,--UG%"E.[R68 
@>071$!8_8LV.J.F'>.,VY$/B>.35<K5N(@()T-Y93XP 
@(RQI]0K6\ C#F%EN(C2-*\WY:*/<<*&+J?%V51CAN60 
@ESSTK5:<!N](S,K70UPJ== 4<M))4L-7PA^5X!&?/-P 
@ &! TLZ$G4W?V#Z5WU82]BJ3_ZELI9X@52?2.@!<6'< 
@;,YMWHI&1M@,=XLZA*\[;URM*XG0,2+&3E^+*90_<6P 
@6.G4?D#S1:03!/2&AO[Y3NF0(*QQ"U';H(._2!-UXM, 
@OQW%Q8>N'%B6KM"<>X>'L^(YT-KN5:)#HI"1ZUIO;HH 
@[W77] 4FU<\.I9=XGX,%H*U$C25X+KB@SN2MZ-54P T 
@2OE0VS-A G#BI-7_)349^S'';4T[MKF31P0CEIF@/%$ 
@ =,A3QP^U\<+<ZKN,,,O711$+^O6;HU%-T^XIQ9;ZHL 
@P;<WF79"P8T&J-1@&,SLI=;@V1=V?K"J%\ ACB5RB3P 
@($MS\O\_MJ--[(792FUX?!A1GYHKDJVL<[0.X;^@#YD 
@_[,BCGAPD*H>O7".O9#U]KX$4H!G5EZ=Y5T3RKQ[UP@ 
@-(\$\=P='3;YH('+L<R8]B_C!-Q5QF_:&5>$?6[P3T< 
@'LL&O .^,\QZVBEWRWT@T,W!O>P1U+RO>;Y]3S0]K)L 
@UJO>:2 G^,1B,4PBC3$G&<*1'0_4Y'K+8J9$"[RO4&L 
@B>P3QNIY18$E?&@[+^--CYZOV[',6RX# /BNP6*T>!, 
@$K6:.F^0^>81V=@%?:S(COY'57=%(ZQTMA4@$O_K23  
@JVG@DC%72Z)8-& EN.OYSU 4>CU]+R.K+CQ+C, %Q>@ 
@*;)V0&!$XEW!3U_L[(W7F+5@;Z/,.&ST/IX^W?)I7JP 
@.V(R!_$.KU8'+0!$]T-M/PN0SLN O$<SD%VD_4. EF4 
@$BD[PP;TG_WNH@=&,#:&BKO-F*HU(("4Q%=HA[%3V!4 
@M<L*9I"HQ5I71*4MHU%#K/AG[AXR^!_ST//#]C=&'0D 
@T>#[2\+RUT=<Y0C*"P70(H"U4<,5DP!K>7W3DL+D?]P 
@B8H0/EV=^[MOQ*2U9!-'V;OZM:#>J\9MU7I8"9E64"( 
@N)T4'&98)C):NK[*D5QXGH92M-EKWY-,SMO5D##1GG@ 
@]W8"C=S2,FD$13_WZJLH=&.R>CKI@"XZ8X<U*>]JH_L 
@7$"X+H-=PIGG<I)OV>]7R&4="77I\4G^B\\)HT//J]\ 
@(L(>NP:4".*TCA-;J+J,;;4%%PVL^-G<V034?%_^<90 
@UM!(2EU ,/A^^CX&%:CO@3;<3&$.R* =QD!=1:#E_%8 
@J1(K^&T6ZX]C3>R7 :/2\RS&;%,M$P)"S3+.TX,0-DL 
@@F99WLI<]8F(H@\(Q<(48AP&[W8^'$2KTOW' 8)[O40 
@F9P]J+S*+EQ+(,5.H[)8BJZ?-/5+ 81RNJ]#F3'LWOX 
@J65E;+L=;';JUU?:I?%[OD>M9%DTEB9K(][D+,T^O58 
@9 [RK!V?%M;-[:,:AY;5<A_.DVV^:!][P:/PJ9E3 RT 
@\3@QO#L;?#FZ(0[_C"+7WDI3%NVP/B"R9E[PWC7A404 
@.(OSG-5>4<8%X^^<;\CS3A61L#^^JHL%3._Q?TBALJ\ 
@<8QWF$-"5SP?+J0H!./2K5\T,6TV2-!T1<5VY)ZC%/4 
@SL*X=3JRYP)0+/L<;!XJ=\1+$0&Z)+X'O+-Y_H)Y:9\ 
@/@"3W&522AYXM48-UN_<PYT[A7F6B[7R'MK3&>/*CP< 
@X5;HUC85QL[N.<Y?W)BTGJW1X*0JAD@5*S[&^$S>,64 
@X8E0 Z:R$8R\OW[I#UCR,8JF@&\&?[#,_T$P8Q:C"/T 
@7S)LA#!*[_6X@?J@#Y!$VKV$.>K&(?-I+Y-U*H'U.+P 
@B;["TN4'TY,";,XCX!_18E/QD\H5EA+HW7,*,W$OK@L 
@ .5Z \%C']R*9)SF;>)%Z34G\^(/;!L7'?8')XH\U9@ 
@Q8TZ"VB1HN_X;1/6TU%+^;U<JY:Z/V\4/0+GAP&Y8E@ 
@"W@B9\;> ,*Q0R@)"UPS"B%_N+_G67U5#K&K'.U8Q/X 
@B$XH*1"XT?>NG"T+3\R>8Z$0 "#F.T\YHMTKCB$&_[, 
@8 &IX.!D[BFS;"6%_.5  ?M^Z6U39E_5]^IO\2Z?=L$ 
@=RCP$R?*'XF,I_[7?;^1=F*:^3H!>R1MH50NF"#TWU0 
@%"4&"KM T@!\(F[U?.>:6MDF!+.I#^!(5@U-SSB&W$T 
@]D(WP<\,W>O6PJF+"-T^2[Q 53Q:!I L!4C97\]ESSP 
@74<5; N.ZP7Q]EQ;Q&U]@YCC+60W98L6@IZ>I2_(A#4 
@4#"\ GF!^F(Q]N3T0%1DQ4T?9Q;UDH#[N4Q,[S*[Q:L 
@]#6JQ7PK0F" "IMVNQG)2G9V^%FJ6O'=JBF1&&W1\I$ 
@:[0"[&9SZK&0VLB8.6=.]SBEE\7PDV"7VR I3NBZ=S$ 
@KAFU18ZQ]8A81SD$]1?O.>+6>E0+KDFNZW"L_J^('?( 
@4_O+F@L#OZ4P^.IU#PF^BL !AI.VZY5RJ=Q&M.57#?T 
@24+N:122BIL$C/D'?\!<=$)9>HO84V("*8$!-=L8Z"P 
@>-"17!PK9,T<\P"7^.GMI9:Q<+L _P!&_!WH$=&_HM@ 
@&]II*<$T@5T_5!P66BL3FCBRVFT7[,(4\>L\B6,.\P  
@Q[5_NQC+93T26:-_P5HF6[8&4G9%/5D*+7DPI@=-_2H 
@^/P/83\0VR2FGL B"4.E\&'?PWRU8^R%@E-^$[C67S$ 
@O]'7?0+&S3<['CDCW(@(XU4]D1<91[WR(V"1!1'AEL0 
@3YP$&ZZ(6-@0R %D<HB!,1WTS*TZ; WQ;(^GZSI(]ZT 
@;5@NY@8_SK(,CQ9'<IK L6Y%^KLT>S#F&"%5BRXJ^@T 
@!<J W/Y'UP-O%T/ZM,N"B':W[[ **P'GNO Z 3A"%2< 
@73Q9V7RNK9\&_AIX/#M;SN3(-:!$2U]:2"_D8+ SE[$ 
@[:$O8'\Z74IA0P@:X31#3<WZD3WJ"N:<J-N-FS7C '\ 
@(/]"</77+=A)6)VK;-RAA05.VYS*2^A"%W]PT]2^3A@ 
@J983-[Q_D.S5$@EPV%(S'(X ^I(8T,'5L?J[0ZBZV^4 
@.E%!  8!.*XF\E/;EL6#1HC.F8)WX-[]8],^^RGW4(X 
@#+5"'J!71< ##M5!]5NB=IE*@J.9FJ$NG<M@O5Q+\9P 
@R*,RND[V1.ZOXE-"^'[10AW+9V4 E!/0K=5DY2/J)4D 
@GNS*)?-?06# M^Q(F18H2-GK5_'9Q%$)6(38RW?\18, 
@3K7VECRF<_8"*C/JO%)(<VIZ^A3 E%3WV_X*L@&I7$$ 
@1(-/KM6F<>(K=7Y">=^@E'VW-37)KTOF?W!XH1US,UD 
@^LK:X!R?@@D.D* B_:%4HJQ@?.A,407H4"Z:\_L#[+4 
@^YSB2KX_]'G&\=QI]SPZ[+B?E947'"T.X)/!3&G31RH 
@'L/#TJ0VTP(I#AH8+\5B\$V=D5+R+TY[SP!>-TMM@E4 
@9YP=\+5SU#N6SNO-I%%)M3HA1=Z0T$-M,Y\8;G[NB!4 
@U)ZKS8(#$B[,,OM)(*]8.WE6O?!8;FR'<9<@"&&MXJ0 
@[T[8B.6NSW!S3I*<CRDV3RQ0D!U34^)Z%P)\^!Y*C)8 
@4MJ7##<L\LIA5..G(2==@B8M#JV*#GD6B[8ATU]PZL( 
@&2LRX-]>IZPR%&VW\[+CB9QXL!I3B/WE(2H^$0>!4%< 
@*"\V"T[O;O\0^^($"E;[-2\?"])P[R/WQ<Q?[],U3D( 
@ QT5'#V0L)B!+\"UFZP^7M POU%I8?03 )VE54+19^X 
@:]AQ");QGI'D]_&>(6K\#>&JY2_6A<(]YWD2/4BO @4 
@L4"@7ZIVBM4,+QJ1Z"A_%B%C_KY@:SDZK@=SS_-WT!L 
@1& XSF&0GZ]U 1JUJF$AK1Y\Q BT9M5P;T&]26W!/$T 
@Q1B*!A&/*#M_F&KQ&D*[ 15V4A1SU(-@(CS) 1<?T"T 
@5R*W@W6R=P4)<?HOV NR WQA_.&E+,9S C(0L:2J*9@ 
@O'9\T)[T7D*>HX&CJ_8@5CC"1/HM&ZO:#F)RXZ'L6"\ 
@7]2N&G]6H,^E:BFZ9+C6Y#WY@ZW".2WQ@&#S<Z$T"[8 
@@#4#':#A7*#+6%[U$>_0M6OI#-S:0"Y_:2[ZZ[%LZ1$ 
@VFZ,0W<KR'"4DDWS.)PD!VD*F!@)^S7F-X.YD13/B20 
@,X <X:U-RYVE-OB1: J*^]D0[4%BNR] 47T 4DV]'#X 
@ML/_N0K-#@UR#(&F9;Z5RWFVM&U]YWBN<Z=\HJRL&QD 
@1U!FH\VK/GWG,VZ^"TNBMTJ;@]B3)AS6L](.(C-N#Q0 
@(.%0>?1\^;YY&*U5W'Z2G)?4#46C600ED>SU[\[$^14 
@14):A;0HF L(R_*N@DDB9L<_GH!J[0K0*@!SU(->M88 
@;-H;(G$;Q"1+OZ6YT/0%;\L&=,*] >GVW/N9SAI7Q>@ 
@KKPZ,5O]EY!LNCZKF#?(PEUNQZOH'*&AH-,,V+LC:NL 
@FX3/2^WJZ\<(/3EH[KJ/NRU 1@RZ7"%P7T"UZ(SG$5D 
@MDQMF"'>UO7_#6B/G'AQM3*',ZZD%%@)9!4,I8LSI=P 
@GL7XO@&V+6JB3 9*D?L+&#*.0%CTI@C)A9KUL*%@JY8 
@\PG,M)0 JIZ@JXRDOA2LKYKGG@RI-LF :9&[I98H_0\ 
@U?XT+\Y?6Q9C G:[DPD(OH9(#'[R.(PU+#P538EHC < 
@N>IQ<5[=[89P23;G,9KW?"$\[,Y@=IX!<H?^NUP@VT0 
@UP_VN&?V1%8#C<VI4"U2V!<W9U (,G9PZR&EP\-.HML 
@<#0 D:^?<ZLF+=\VLXPENK/I4"BICP0'/'M@ /R'EK< 
@@0!Z#SP9L@%NL^%(A6G5,L27A]*PY@$[3\!.3/=@BX0 
@QNBE>*B]0I,"\9EE:DGU#OD&U?'74;;-K S.Z3P$=*L 
@ALK7>@ZI&MY[=V^0F([D>M2H>50 VD'(E9$ANYWFW^T 
@LZ+7;?6]-"3':NR::H>6_#>NV,T+Z0!2%I-SGD>'Z2D 
@D2:AET92^N9[.,P;8!""4 Y0NP]U;#S/4*<+CB&]F;X 
@>ZCL]S!O Q GV6SH P&3AZ3N8=N-=/*^P[?IWOFYF#( 
@92[0?^@ #;C#!]4IERI8S!.#X2XP*R^!KR;QEM%2&'0 
@D;E.78D:^<6"]9"]+*D8&^IZM[;4(_HXC^+;J]I*AXH 
@!.UYX5I', 2>P,C@<YD?LX]QB>$4YMOBA-#:5P:FZ&8 
@ZL\2_YW#)F[@;\B_* ]SF6XP)@WFL*]W+0)WI)-#1.$ 
@39O_9)4)7Q%MMN1RJS[;B5UO\!IGWMTW&YS1.C7?^$X 
@1QJ8)^'I;>0J;,6HUU>W0$90EC5J,]VM"8<"2T?2N!L 
@TOS>7*"1W9V"_.J_O=J)>V&%@JXSN':I_]T 3XY=[<\ 
@MEPN?!\;K@KZY4V ;)Z8$X8L=,KDC,V:K6DI8]?6I4T 
@KGH]TL_;6@PMPN -/MG$VX!G. &'&-GTUWA(2D_&C4L 
@)@FQ_#1I\;#74Z1^:BV$JS;1[=8&:!!DZ@,U'HS-FP( 
@(C>CH;*L8T'?KQADQE#CY)> =^GA-,U;_HC^+@3G/2P 
@;E,[CA]>COD<)*AT8VH'US]4"F^6<;1/ ]K+I[3!4Y, 
@.&!-XL^I9A$N"+M)K+GRZ(ON!K\N?V!2'5K@@U<,CLL 
@42HGB^P 7&J\WMJW_NXWY[1E(.8I"9Z!YKO6SA!&H_  
@/O+8C^<*JJ$4]!;_/LL>B1"F8,*'[K':YXP=;61@M-X 
@I;._)IVJ/S'4('UL;U$;16F#* 4_XBK-,,?/MA/R?>\ 
@**RGTOKE,_[X[EW 8,YD^89W+_CAZ0-ZTYDYCY9Q"/4 
@X23 FA[W?C.D+GD!2_]#7;6$D(>,)[+SG/@6\/"&HO@ 
@H3A!E@T5,)X,Q)G)W.X&)G$_ZC#7@C"*0._XUIRG>W4 
@-1(P^4M 2^(*VO]!UH+N.U!#3V (WI-9;26CW=)M/8X 
@#E1J OOEDNR?_#H+\$) @+ 'F;N?^SC/R6K=YU6+S7T 
@IQ'L:2[:MP)R"N(:]10;]HID"T=J,=*K-U  0-!?S[( 
@R-Z)];K1*WX:Y,P&?32'^EO$(0;"P+B(A"7U!P@_<V@ 
@F^N@_YK"<./?FM;#07QZ5O4J[U?5!1$\:]\&A1T*XK, 
@5CHJ-2,95_;[R3Y]O9H NG">NQD+6SLGFF8W>J/T19< 
@4"ZC8M3 K.F3G29UI\+90):YGZ+A4)1SN\Z)F];J^P@ 
@-!E*GB0%]/TM@0(-=TO/?9IZE5WRX*^+M&50SY*,E2X 
@.W![GRTS&!#DI8H34,3N4$[8)[I"PPE(1!P[ K8*LE  
@JD66YDZ>HWII1AFV#O_1U/\R,BDP^4.([%,YNG%5=*D 
@3&-ZS>K7=N47MK$5!Z#4<\:ZYZ4>MV2;[BKQR4_11!( 
@ZOLMV8$_<^-&++ X:(!<5=/T1]@EDU:,R@L*Y]:CBR4 
@ CP#BL[]F:NM@UU\G807ZY[/ /6W=''AJ61EUDWXSU( 
@CD"S)XS.:/%@8SVM3N%K8IX]PE)O>5*BI'H1=[J-%"  
@S?;T(2Z59]:S/+:ADV9U/KG^H9).*FZW9.;8";98)U  
@G*F@?AV*.%>FL1QV6/@J=RK1H2!HYWP_7!!C@ZA]T[L 
@5:Y3ZW5O7GAUQ8P/0G.=+-;5\B9^E$9IAIM<KN?)P]X 
@AIG2\<M2E$!MF/Q'L8!XQFXW:U7T-/QNB/S-K(58!=\ 
@0JWKZ\;I/_\=N729H3=#BA_6!8)I-9 [R'38][CM"G, 
@%(;L0G*SM[=>AW+7TQ81KT-<$_R>FL,W!53DJRL.F%X 
@8C[6#%X,QUSKGNZS2)1N7H5&8)DI4L\1N.]7ZN*: ?4 
@3QSA90$XZ !]-RCS=-Q(H<M<#+8T&MK8L@XOM'#*^E  
@P?CU2Y.J.*6B"@,5X//@8?'1>:_SZ2A*IG*Y'S[C)24 
@F1VX]=A>YWKE[Y:!JZ\ ]-AH#G37C7S9]O=HXP08M%4 
@1J.IT!_5&/ CJMME2_YEZCD+W?*?!.'35&5@UO-D(N$ 
@0*32UY.G):1<;?& >,V9>%455/[^(X5OH/B?)Z1)H#( 
@BPF9R3 E;.*^9P?]F-GZ%FJ[@'20+.&TI>IV+W[-_"( 
@T?@8RC*UGIML47=MB[(]#LE% $UJF&<.TCOHMFWQ!X, 
@1TC0O0II%)#0TBZBLJ8)CS" H&$<\^3HQ-A__<H![TD 
@S;+CXLQ7S*L[1@U[J?0?(:?V2O[>QUC:.TG5ZBLT;]( 
@5LRH'<H>U$^<BJ\6&TJ5GU<SQYWSOSB[-K^<\+6>P-4 
@#DAS@C;;)UMQ@NMJ,$B,LYWZA:MF^B:T/SJ1YZ+%<18 
@RZ(PP;=Y#PIM(T4+SKCY*GR%91VKBD&4HXZ\OINTW<, 
@*GA8QQI,JL]"B.V*(5J?H8&'<XMGO,,J%[Z-HP7V\(( 
@A[&F;Z)'G@82[V!\&F[7+ZAR597JI88EYD.> <#[<&P 
@%*E(K 2T8T^TEG"FUAA>8V#KA0!/GPX4>JKL06IS3DT 
@NBNTSB3M?WQ-LO9TBPU]=%<3(R*]@/9SL3=M[@"?BI< 
@POU/R[.3<LYYJ<(Q^:)]@="WU(ZF98-!M?!0.Y<=[=X 
@&Y+?R<0GV9L1*-+<P*P9CCLOQI2LZ[&X),_VS23@D_X 
@OND*]0XNB+L#9EDG1$"O]\0%=O"LTG^!9*C2,0LEMZ4 
@U\)H&+EIY&?0I4.-ZF<24J;3C5>:$6.CAY6RCR4]%-, 
@6;68Q!%_ 5%@B'QG 1[PGPB"VI]"K!2'5EI*LJ8E_!D 
@9/\69F@%Q?O#3E>K<?+(>I60(7=F9"0PN2_#W:#$!-( 
@V]';EA]&W:H.<A$O)X.F>%_K]IBQP.L$?(Y%V186*OH 
@QP0(Z (._>$>GG"C<,GUBR,R@GKGFIQU(F0I3;+SXC< 
@8EI?;!GUH!][5$]N1V<AON069^FZJN%CRL(KG#>:N?4 
@B@*<EF'PCP]J[%=^:A;>SKOYGVY<A!RC=Y7%X&LM=S\ 
@!&<KD]T^]$'GH31>>K=HU#@.BQW%>T$#?31!7+]N\9< 
@/@I(,4'-%=FTE>D:LGG2_&E(D38*GP'33XV?:YAP@ , 
@RV<!GPF8(0$54Z;PYK3>N\CGB'X[BIT3_B+U>EVANL< 
@.@EVE<R3P_,-JFRQN6&2GFA]<V-@\-0G(!PE%F29%ML 
@>PTK'HQRUR2I2UT7M0>#4YD2_\Q]/EHR;[TQEYA?\SH 
@<32CD=B-N;(4#XOESP EE&\]5D&:P85&*D>ES5<U'24 
@R_]O*-K()-AUG&4/T;Z$GX03V@21G3YH8@\'EISX8EH 
@$C_,1:58(.D!G4A8G@\0A7Q2R84Q\-)RLZG5HJ"#DG4 
@,P]@B2+DJ:<]<3TIIEADS4$@'!<QCYI69CU24YP[S(  
@7V"%U[@G;R\!9B+%<; YBRL$8R@P!NSPOU?Y8[W0NR\ 
@!\71HER(V,3.&Y0T8H7O4WU)LE??0!92,F>0+AOZ[N\ 
@OMX.^ R*_?J'SN1Y#+MD)ITKQYS=5 4SV:M%JC[&L"< 
@N4M^ L^#4M;7DV+JJ"4)\-J.B;B8#G4CNNUBRW<@A P 
@5^6/%U\S 3 -?VL+5;_O ?*%(\RJ1AU)><>GKPEH\/H 
@L62EWOBUA'QW-DY@E<.6\65PV7A(\%NSLETO;0NP!X$ 
@[B[[TP? A0M51ZC6W!B3^LA3^_,SPT=T#WN25RPOHV8 
@ SOMXBSY$B:='>@R3;TT+PP4I33'JI 3>$[10B1[0;8 
@>I-'N$G-W P_<M2H2V2T5 X,7K!B2RO^YK:2C&?6.8\ 
@))^50#FAE_&^U+W7;E\J"M""BW23/_,5*ZRY@/B7G'P 
@I_IHLPQ"UQD8O/VDM\ 2XG5-*]\9@BT5X;M5$%]P86T 
@QT8JL%^:<UVO)NCNB3Q73+8-B(S- N6$_=W1>A-/\!@ 
@5I[?;;AG5=Q6K=+JZ9Z*DEXQ?FPB9B6$VHENGKBO" H 
@WM:<X@"RO\+!&15G@"?B<J3+"U8Q7$B#<K2;_OI;O^$ 
@/8E0"V]\(Y^81FI56U!P[NS[/V=2D\K?GO$19</-,:( 
@'ESZ+C)-O:>PFP9+P_O1#P='G,]=-[F?-YZ#R,]S=7P 
@O%^_ZX8'5= )T-1P-0BUUBW5]K<R!(!ONS@?X/T)VHD 
@;OB?]%_X 14K3R,3,P%N5Z4O.JX_.%= A]I,F]?>&Q( 
@:"TAIO? *DT?&PHCW^I^=O]UU-:Q6 H'%/V J0E5\_< 
@K57K]T.O2HK_G-Q99S))A^WX<YOO;O.XDHJARN"1EMD 
@,\ *S:!2>'K:9!A72*HI/3T;X1I^3"%P(2)NSW)4+NT 
@3?=Z>Q3T:FI&O3#/+'):$@09R5B.D>UC3V_%:0OBLLH 
@A .R$_C?%;3BKB"7.TMW."6/[L^7OY#K31$I!KJ A_@ 
@54TWFD[%/?]+!LC=AAW>U9T9V%FS[JJ"4TR7B!\;W4L 
@5(:2KG6D89TANK%% P]!_QAA+;#=!+YZ58=7#EAQ)&L 
@*G8S,QMNQM*NI6V9M"*0W%\8:(,74R4\:NI:(Z6DB7H 
@7:KBP&"Z,-$\5?8=EC8P!GQ%N;>F-D.Q%Z]"/3/%,GL 
@UYI<F1J#5#QET)P42C<+W:L&N)):Z0V,V>'FB%)L#(  
@*PYFTW5,XSL@-V\I$2MXG!.Q$2;M=2^?8GN9JT&1_QD 
@0OP<['I4 Z%O1ES"O)22EX\)RF#TPMTL/89@\@/% C( 
@,RW8[U#VJK!^2+%#W=WYW5MJ_:XC;'FR8?4Y-MXD;F( 
@%:.8U>EB"MS;3[E$-I=.W9P;@,7I_I]BF*)Q9(\#OBH 
@-*Z.>/T^?*_S!XS=FUD2A2M!P'S&VWID5OF'7=7YF/@ 
@0X2/K9)&7VV787$5C8X?$%M0$A29^,O\$=![4HMUSLH 
@-=>3 I1K!U[+GSJ=-[V O&J;LP#>\SVV5MP*1<>N< L 
@L\NBQ9I1!AQ%!)KXM- ^2B.=#.X$? )1QY]!EAC=D&, 
@]M^4K0!]]/36\+)JURT&JH6YUS1S()U\G%*".!*;^T  
@"U0 A"Y<1F\7IE/FU%:&>M<5XS:O$FM8CQ?+7YAD.D@ 
@\)/5O*/N]I Q @JKXB@=Y95JE#W$!O\5= X.8BW@">, 
@L5EU$_WGOUL%\/+%T L"#KA(A2FM=3QXK^8R2=57II( 
@_D6G7M0L.5>@H9W[5)A<+2I,3"[L^G<.V+F=6!"^56L 
@8;->?SQC4$F\@&]^T=WZH?LIGPJ@L2;&@68K1^'282L 
@'*/E0,E3_88:G9TIAAN;6_D\:_^D"-A+3 4R1>;:C3X 
@ ;MM)3*9U__.VO2=H*#8*1\RJ[:^Z K_"875!V$*%F  
@L//1E2"SO->1,^6:>C\S?QPZR9.'#B$ZNE2.O"_^1+8 
@D\06E&1IZ1YRC!-&-W6/2(=H::*QK.T-(&X-%)^4G$  
@UX!F1 7<#Z:%&=_P$-3#\,!):*@ T@6^?E?E[-UI@>H 
@.SI[G=$1H^K@V?V3O1N-"3F-#,$,BOULK!*4\U1K$<, 
@JV]X#QN:9A61NMK>![Y@T:M=@IHU#2/CU,<(Z@MMI"L 
@_\@PY/4K-8#7+TJFIY!Y@3ZH^E7]U&U>\6(EW6U%@,X 
@B#7-V9ETZ@@H@H'FT?B_[QQ[':O]!+CYGRH(&/B]'JP 
@SPT)]LD(3HPH##:\F2LKRYO>75G6T82L5ER>I3(7,KD 
@N)4UV50KVIT&W##[+XYSD>,9\P _:K7V*>]QZ6A,D4H 
@KNJ3=6JH;FHAQZO\_:V.?Y_?C[S">'%>\'U(ZRL C74 
@G0_*4E#!C:]4Y4EC-$9G L$)0",2/ 5SWOZ,LD2I&Y  
@!28O+I:D:A7P'ZDI[%F<OA3/Y;'21$M$,Q@\-;/T7"L 
@BU3DRV7,&T9O.UQ$P /+-P1;N&_YY+EJ66Y)92UN5G, 
@I"_X+_L[RSX@4_61Q\9J]\1/'1-C,2C[3H6&#Q_UM;$ 
@L?P+C J=>A<@SW5$:ES\X0 Z#HYCVGH3F,5E#26NQ?@ 
@  * )$5CQY*?T?]G_4ZB:ZK]<IM%&,&P5(],3BZQ"]T 
@1S;I3*(P%W";(+E&NCE;(>I5V0D4E>]0# .TLYJS0S  
@1U1.-TU3P8\%@%>;7]MPN!:2&US:>%5'4\'.']XL4XL 
@UBT4!*CC%R3FY#J,Y+2I->% Z72^9IN#*SMH'3A58\8 
@T5P%O/^S,S^RVOS/$J"H).[C65M(A.-[.:Q^'7<<A<0 
@3TA=3)9=SN--J4F]U5GFUXK?6J&T'$U>W5DBG/C=\2, 
@&[ 7$H(&8[OD\=32@2?M)U=)Z3GK#S-6,8&6_%TU^W, 
@<P>WK[3?GGC<S0#MB6CCP+_"M$Y:V9%-+MYYDVQ*<+@ 
@M')HT =2X  EM53C[ABS'5_!1&]UAYC\!=!'7"D=7A0 
@*=H6M6<1:VJX5VGV5(*^@W6_.*.ARPPPPS'5^/R8XUX 
@JWK#%USV.U(=71H )D(YVUXXF@=#%U*O5#W 4![/&88 
@WF7XZ&B/)^"NIVV)?U;6,CK:PN>SUYGM?RG(T:XMX$8 
@+KJ_D^@O3M%S5P9%'"SFZCZ"MN/Q.=\K_ NVIB1G?\  
@\O>FSZ!"V): 1)2EG7UE@LM'(C3$XJ24(89 G9ANV8< 
@3_@&6UHL'R];'&D1:(M<#.0Q1S^=G)R=K^>#Q>BX#/\ 
@1];GT(53V(V!D Y"1):SND4I^,RSG8IA.$DI>N/5$$D 
@8"H.0 V5V!?#37S=X4:).[RQKY>]_K[>XMW-,W5%<O0 
@S';/8T4-2ENW5WZ9.7'D".0?0;CSGF4UA,MME:-"0(, 
@F9@N)AL$)ZN7!D,;3RA^TY@^B -G5-#0J&-PI'(45 8 
@%@Y\FC1L2[\'F\FUJ9"?U=#C.@'WGND9[]LJ1.HX<74 
@T 8IG(+F)K9_)4E75SOYKDK6=3D_AT5#HTU#X(F@D>$ 
@^Y>['YSR6G,8$DOU1-IU\LWU_4HYT_?<1PK33[)HCQ\ 
@%4\% W*C>*T%HKC<_6S%J*4C#Z=1CK^3A@CJBO>YN*T 
@+DPDV]P!N=^75*&EM&=(V=O#R_O?V_KC&;_N)Q8B0HL 
@;!?(4=UQ&093#]O&,GSF:[/-"U=MCOVITDR,<JU'\-T 
@*8.M'>+!J;+^X>;)=YJ**B2?93DG<I BET-MGG;I6Z\ 
@?7"^DU6&KTV=;7J/'PL!BFYYF_!,.'-XBI>&D0,OA+X 
@EP3;O'VOD$POH?L3VE9-US.9?C!76OC\8EM;E MHD.L 
@5S4I=.%-@$A!W-R)4=@!. XP@DTXRE2/1P8AW"0+P_< 
@E@0T==1K/F]W5FZAC@;^-QYULN7@[L !>G&O ]Z9CY< 
@*8>62WW8R9]G1PGTIE _*DLMI=0IK>TCF*D*;._YU9( 
@6Q?CZM0+#*O[8&-K*F*4TJ@9E,EH)NV_2"C8C+#A[SH 
@D,/,.D&]0T"[3OJ-+_.0\7%6DU,A[7YKS8^?=:3-. 8 
@<507V00G*6&L2%I,Y3[>'!,&[!CYN<^?OH*!J&J?.E8 
@HX'IY @IN6$5C1<;?'Y=6@7A:SF@W<)3[&X;@TE())$ 
@&#-B!_)(KU8"9%\T1"&UR$[;##)B@B\;"?G%9X?&KSX 
@Y;%P#O0TQ%]ZK=R'SBP-_3_I:KH7(MS"@4I@XOHXXOX 
@]\#=]6E^T9"Q:PMB(%Y<KA]&1V/<M;^OOX5 L9^B:K8 
@9MF1NEJN2MPK?)",S6_:>G^=_\O&FE_.@76Z#@/\<Q\ 
@XW M O$U89</24$;E>EER29SH%,9(O=ROQJ&FQ%Q_NP 
@V<TB6B6J#C\54P#"KV4SSM&+-'%"P8)J[!A";J)S?]< 
@(-Y[\G1]W0R6WRB)6Q7U+9PIE!I_@V3J(R6N<\[9:<( 
@>ED;6P_RDNU)-36I_=YKW?J&'AX?%+^4(+71.E&.Q@$ 
@J7Z+I-RK$8=/0$)K)?$UXE.+NH*L5& R7(8ZF]^Y\E, 
@\\&50<*[/;7AO0TWH-[RN>_$MY+UQ;KA+J=E:RJ@"D$ 
@<W9F8.Y!$J$L^1<)#U<A8Y?E^K)$,:Q;IS?18BHKED$ 
@[6[PLP^[ 2=2;O?S=9^58)&;M;0]WL;D$%MK3%)$V_D 
@&J#O@27WT*]=BF[""NRMR>S%6>"% !P.2SB(IC%NZ_4 
@JTU$A)>)[$OF5D1;N4\($F/Z()7A,N5I@5*7ED*C+L0 
@&[P?08'5F5]&O0?,+=$[XX@P' Y9%[N_@,I/4!J-)5( 
@N^FB7&).W_[STW4.0GJXU"E.<7A-M50-_H],3\6 WUD 
@+(1*99L"DRZ5;.5IIZQN6Q],5OWDO=2,2YVG0M:6Z;L 
@8[*W<\@!_>;(D;'H*$4^N7ZS*R--EQK@WNX>[L28*4  
@YLA8(O^K8"70A/WF*B\,?V_+*=C[,AF>_8&5[D6H(1, 
@7MV<L$([!!'/9E;I+.N(&M#_:7\X((/%?8._-D:Q0S  
@+0.Z.$N&R]E\\F72'&BYV:.)9*U<XS2^#+"K:_-9<M, 
@#Q<<S='&$G=$WGM]RZ Q=2( WE@G& <S'!=GK,L";Z, 
@D3>H4JA<:-31[_:NZ/CMSE+\_*\;<^CQSKHBFH]":W0 
@UIVT'H\FE1ZQY[HI[@3]KZ"B!?[U+(#R(Z(C_4$K(H( 
@8I@0$71Q19U>>RUI5X]>E@^/O]#PF'7,-.%LHHJE4FT 
@N UO\J"PB0!?="K,;]&70?UQ42N8,4Q7&#1GQXPV&/< 
@S5'BIWN5(PO&P0I#<L$A_E\<>.6Y1J#V]>WE5;.)76X 
@8W5-?ZX:FU=8N40N@O@D)%[ C""-RZ,97<Y6.WY_Z,X 
@ 3B@%6^"5XZ/WRF_ 4GG :2\0+7^]TWSV^\41@:GHC@ 
@ !#RC%YQ,_D&AL6[Y5:V /*C6=7CVJ"FI1LR_+>JL)L 
@UC.,]$+=-%;AUEM3<O]_L'/E=RDAFQ1UZNE7%=*'K(D 
@-IU:#\A7M5@#C[4:D9H0^SDKW"(7+OS$ #Y*E>BA$$T 
0(!9L^^/E%Z+X:B)L'(/[B0  
0#J.F2;U8ND(#S6+N,ZRSSP  
`pragma protect end_protected
