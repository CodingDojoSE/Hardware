// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HKD4"@U4]0:HOD+^W=+UYL7<H8YA9[E7+4R.8D>XXB>V?'2[Z/G&A?P  
H^H+ZGSR6?.XDV9^^7H&>\7#'PD!WW\$HL%U/Z*&9MT'T>K+\V9&)H0  
HE%WJG"& [JT./TE[?2H^.6^Q76X@/LBA[6WM\AOXL"W,]XA%QZ!YU   
H%7,C<J(8H^X8RI^_V,D>5TH*7!H\N(H$V6'%CO=%LJA,7#;M*8SBG@  
H5$+&<+.49+1IJ6_4%3Z?P=K$V8-^RFBI@J<"2F5V#XOWZ12VB,FJ\0  
`pragma protect encoding=(enctype="uuencode",bytes=5952        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@#Z4N[=456)-ZJ(9IU=NH@*>7 V>!HSSOEM+H9C"D&[0 
@R[9^VVV\A3+]@_##/O;0XN1CUO.T/)XYTH#RAY3O.!X 
@?YO'.NZS;ZVX\QZON&&Z*6:&Y2=P9>G$*ID?"EF#TM4 
@L1T(PU%DTPAG?VL]W0JMK7,Z+]X8_>?;B& ""*)\QBP 
@H/AE%';?"JWA/YK_I.4^% H'/PVTRJ2+!W3]SEF4:W, 
@5J#>13-!]2 RK#!7X G:]^4_W".#N=-\/>$%#X9"F9\ 
@P5WSO6@E-<R9MS0)>.<@F6%>ZZC%<?_)S ?PTG/5#G$ 
@2&%\C\+K[6G!*56S,)[1P^*#=<\:N3U'LG)^2\?JG88 
@AI7)[EHCKVP^Q@?PBU-B?>-TK55%IZZ.:81.<N96\H8 
@:\CUE9AB%Q47?TWG:GYP"5 W%H]G2_&GT"FJ+G)[\0@ 
@AS:W$QETZO@^$LZ;R6BWXW*V+%Z=?E%4(O<$\NHN"F, 
@SB!1MF:73;NP&%/\%GCO5U+"I+V(F8&&CN''&3Z-AUH 
@.\X52)[Y4[.*2]'.\S4AS/7_Y2E%(=G!7#6.*PX+LR, 
@Y'9:D.E$2RL<[.!$16E*87<'=;Z1MG^@Q[N]+>[8@ML 
@G%V'A%O)7M!75"V^)V UY!F]9?$& %;"U_*C_L4=-0H 
@::)U;9G8IS_5$D9VMOX:3\:XN?V]7:8?"+27NG>'^O0 
@%*\B(6<^<,W,KN'+C&LTD\?<^<$._,JR&-RFG$&Q$HL 
@\^]+@.%Q%G?,88DGY56PN&XMR5-Q *V^%R4RJ_TOQJL 
@O;;!S-PN#)-I2X8QDA[5"C"LY5&,0D2VEKVU2]I(=<\ 
@8<"5"(G_A$>]Z)NB_8]6ZWOR)!\,<Y>8YGE[,U!J9R@ 
@80LZPC)U1W-&"ZR*PT ;-=';T'8#VCHB4SS+%;5W)X4 
@HFWVZFZ,@5Y6..2@C@8J9V-![O_ZI^NN(.EXY;FACK< 
@"!GBX P=?I;,5PN16V%9^.3,J_5(-WN20,,'$IL:65H 
@+'@8PRCNO0V.))HQ_5_MM1KK>MEF2J]V/PD(F=$-*U@ 
@._S[=)<&FD;L4=\J#3)8P?5+]YU_R]=II7@(;WE_@S( 
@ @A(,0C92XZH_IGI<>,SXGHT$O043K@'V6:*:V?D(WP 
@A2?PG@,3MJ$)@&;WH*QJRDA",[B)6N3/7I45<1X9?<  
@LKYC@(@=K#)0-::.H6ZADS@U$83O^M7<CBKSN^1*6O8 
@!D^1K.)S^!P5"3@RKZ&^2#8[7?()4N43D(BR)3E5(=H 
@ZLNS:J(<K2'L8I-[@N;O+GE96V0FC: 6^_E9:U+#@2@ 
@HP[P"2CD841J5?WIIJ8V":AJ#_OMOV8_U+L4=%D"?4, 
@['=9:_4^88GVE>:AH6\AL*9G(X4$.D/PUGG>6BF[%;P 
@HG$!K^NYOXQX5<)K,[<9T^JNFIHX&'P2[M[$F#/"J8P 
@-1^8K?%X"-^M-V8C>=%\[,<8)GOV)7=B'3^^S51%*C( 
@ANK6*O5\CU%UJ:,#1Z%$ =IVU8Y=OE3K*S(S7H=$C;0 
@9EH*L)D>RM,/W%W4@7@18WFSMZ'BD4GC$Z"@[8/PUQ< 
@LFI"X]N[I5X:S).D[P?J!0VESWX+C(;?FFX4) #@FI, 
@;UD>!T)&+%>OJ)=5RT:MALC$3%79(WN.Z.IY7\A_N&$ 
@[. 1-25)'%SANF-DCG[&! K]8#1]IG'C>+>-L$YIC&P 
@\.@<5>FH4#V0&=]-3IF*Y=GPI_KA:6X-4*/1V-$[NE$ 
@B;'Z.*:.<\J&4_#1W/R';ZFDIZ1K=].]I) _'4HF&CX 
@G2,;B5P+Q8_,;1P4 XL]<4@"BF?%&K\-2!7OSAPQ7T@ 
@OEBHUWMGO2BC+<W8TPO8T]!!XC]/ 6:=4X0BX"#==N0 
@S!G4:(J\R4*]R('2YSW/PY2Z)M[S52Z9![H/GQZ'@"T 
@9$:OXA9W#5QL;.,8@\B3W'3L^QI9#79CWH78TPH( MT 
@RSF!36+-78:EN?)'2GZT<-2&6R5NRD%>E-W]0V+P>HX 
@*D9&KW'(JJ2D^!5/U/<8J[XPE:(,*#@I[*Z$ARFBQS4 
@'J/SU^Q@*8"!%6-PNL$CZ#$C#UKJC%&G0R3B78)^P(0 
@ $*>Q4I1;?]7,5<$[HUD)"Q([SGBL&II%NQTE.WEVVP 
@1L,[/?]-C4C]_VJR04J**]).%H3(BDJ?X,?ET-7U &8 
@F@[NC:P*_KW-[)]434!W*@VC O#>%:_:M[JF[A"+SE@ 
@X1B%)Z+;0)][4QMD(GNA3V@3=TX:D QTVK^';AD'4YT 
@']12T@ J^&2YIVP"5!FR6+M3S+,ESMY'X]@]+UU^@QX 
@M[GD6>S]LHGA_NH!&=,L!\[%RO>"[6..^_12N> 83W, 
@B!MG.L&*3E>3T\QDR1-]"?($?9YU9#%T3,=\$H/]%X< 
@65BU4X;NI?"-3E5B=C[G3?X:2W@SNSYL"][=.MP=C*4 
@V/MT+RC#97+%>06&%,!;>D=DID9]*I  EM'4+^%? X8 
@@M9@HA@V >WKO2RB;@2:Z 2/":03\NWE;FEO X3TF@< 
@XVZZ1RT'KY!_[4OI=,#_YQ/CA,F.!MA10J0B W_2N3( 
@5\U/N[<QNVP-@L^F AF +J(%4"\4^(J$(OZG;/US4WP 
@O1E?=B8H($2&BRK85'733;7JH,F A@B<<FVO\]G.HY( 
@I?X'8YD&PB\7;=4!$#Y08ZOX"JE<#[_'HBS9736 DG\ 
@K_;[9-Y K%,_D)<,XU_:O? F<#]("_3(GV;4QO81GB< 
@?HA%7,E02O,8K]83>*)P[^# 0 Y/:'4UDR=.[SL,9J8 
@7[J+/.G3J#:OOH2_GEW]@ME"'2RN)#@;D3+/@Z\FM=\ 
@+Y!FGW!_O,+8;/^&J+]7%[(>,VFG&\4YWAP E8__NH$ 
@I:0'3*V-8W[_Z.B@9K[4^YI<(<(.2H/GG?-054BI%E4 
@WT%%M_!T96A9\Q=D=7FTDUV V]O+^'..&+?2=I5@*[( 
@09%0Q*J!,RJR"97(?-?=KP85"Y62U9SR^M:FKS+:^0X 
@D,"NBU #W,+=>N&?#<.\TK9*Q$F@NTA:2WH_K,HD[BL 
@]%;:7#K5T@:E_3-M+>7!=(=J>E\>UHRWD*AP\0X3'W\ 
@DOX/=B6 ,[D!C4AQ.1/0DRZ?Q>)7+FQK1+Y?Q6>)_[8 
@7J])R.X^;74\Q>Q4S!(N2Q9#'^WQS*Q2"^9[PX,*Y8\ 
@D5UD'59AC07K=6R8SE-+'A\ N:[X!56X+^<?[KM[4E< 
@%)PO(88#0+@@? I$MUWS2-U78]_['7\;A$A4>.?J]SL 
@>DG>)S]F1R7%K7YO_L>6I[[6=Z //E0 49#=*;,VJ>X 
@K5*27</EK\2U&Y(6F03S#%W<% ^SO._3%QE9:TZK,/4 
@DF?)'4,E_?/M?#VKIF]H/4"_S?6.$ E]HA0\$1\GZL< 
@<GU. N<P#8S_/C')P1P$MAL8; _I^JG2'38);T0O[60 
@+"*?!A8.39,AZ&C.3/MR%]?_I_YM.IOB-EL:AU&!+#8 
@,(H=E "'4[I6B+A3.ML/QOQ2824+.R1I,@T*P@]E^E< 
@<BAB&Q"0J)_.0DI/-27/#,EE@/&FTX#,%O'H6;0EM5T 
@MUYZ9), <@*YT]K#JN*%BQX\9TUFN=M?!FW RUGAIQT 
@WY<D@P!)ENN] <7178?B<(,GR*@41=2!3K'7E8S9@ P 
@'YC"V1@Q\2*C-XJ_:S<=V"L>0LVL';JRZRM=._[MH&H 
@[^'W@KJRZR^:8<)P)+6H(J)(3[](7Z.F\<D+^N&W%:L 
@' ;RI";=L2/(0_>O$.J'GTP_)^7 PDXB.SMJ(XPCT&@ 
@Q17WWL).4Z?"#* >7_73WI'?"LFI)1AH4;'\H=@00V0 
@6!'8RY8?#JAYNY)X?(Z"YZL,@GK34)&(LI*F^EF&26P 
@6M",&<%[9E@-AX_7\NONF38:X^TF94\)ET,DR45:4)P 
@T/MY?^XVD00JSYY)E>5DL8U%9Q3MVAIWB.9.K]]8!1@ 
@)<TE B1'(=N^3N1!=3S,#(!^^/0$!'A[F8L]L*(S#6D 
@BC#D0XP2BZDQK=?!:BZ,DMD6$-NM] #.>DJ'VYU^RO$ 
@]L0?YC,8^H]>"#C<?>;,3Y@,6'$6YZA4M9U)<U_E -, 
@<7W\N'F(M5S,$/7F=.181*4-\')$^JJS K.P]'.MM;X 
@4]1)J#FK)0.RGRY!$'7>8N1*),':J(@/5ONCTSWU,Y( 
@%^QS#M[W.4$^K#H_^?(8.=PMRRJ,/=IEGUT\,=(,&<$ 
@AIOYG,84N&F])H1/XVM;Q'4*T=2JZQ_&*4=#-!:43_T 
@'F2/^UVYY4:!0)88X#'J-7,I??Z)63%/L1FXYS'>PMX 
@O<>)8#FDFEQ4>$$EX7U2C%_R!.RYBVQ_()HRA#VGL9  
@_'Q&6.#E ZH9GQ>B2!%(E$Q:R;]BP.>C[_"\GS:7%;X 
@.51\)F*C(T5;1SV0B\^UVBKEF@ /D.UE^?L$5X3'^C0 
@$AU!UKXV$/^M9(L+O(TH<QKQ4FHE6Y&B?CU'Z_T8IRX 
@%PG*T!,@8LV"^& 5+; T(TG+>^+KV@4"&7L<6F!TQ6X 
@Z*]\:#3<@N>64:LZ7PY6*1$7B-W>PYG@P"8;-ARAFH( 
@1M>^PP4*[W-#U$])U=2R;52W_4"\KN=FO%;.^'#14PT 
@I(,KO67\Q:(SAD$-<=':!]U4RBQ;@_-4PK,(&JGAXK4 
@+<L0)N@ZAA9:L9FD9..08DE#S@_.BUM&<'1O!"&7?*0 
@#M(J@EU!(I?U_;K"FM0(&3T\V:&_ AW]GV8!% H3_C0 
@ASE64]+FVV:(\:.G9=^AQGFU[MY03CTRBC1X[D^G5P  
@9F_\/R:@'LKC*,G"=0[M().!L0<MY5T:.=56L,_35.4 
@?(+!%,>3X9JFV:GR%6L_(B%X07/>B8=AVJ%3"_F!^#, 
@%C#A,)G>"^ W-;[3DJ7G7&DR6BRFN9?M:=J8=D2%50T 
@6):"23[8G @_594KU2S:FP9X3*%/MCC(9<AKT&)3(/, 
@*/$%VZ[OU?$X,;1SQJZ/CWL(F&F[U,9'9'*D*$:XP]X 
@.)ND0@"1>U#QY(UP"MX]7[[T,Y"-2 F-?<I11N0DI1( 
@'EHQ9?W?CBTC3I("KR8VD.<N%.UPN1PI8R%IJOLD6I8 
@,X7!6VO?G#@FTDV?VLP9Z_$[FKJFH'X5TF-A *^@*=$ 
@K^I/9?LBX#G)E9/6]H /VX#*,=#A(.*^!_@*R*(T(,8 
@^N3*R+P9BFF!"\J3%'!'N/M1 UPX3P'$6O8N.)=2DBP 
@IU AB.1Q;6_XD<3D>@A-ZNL[M4RX,?"MIX&ER08%S68 
@)X,% TU77[V* !=HSYW2*>: GBZ^NSD0"7,F9HJW^?0 
@.3W /[OOK][U">T&9)@I&!$3R=?1@<< R<>WO:8S$Q\ 
@6*<"'NZ"<W"S#Y5K*D?M=$4*O2PFU;X,HC;2R\G4_'X 
@'*Y_2^%GJE0%D--J]DKPH#B'9,PR]E@E>Q>UPW2%?ZX 
@J)"1=/M1J[3=1WXH$)23L,-'_3CY"%:0UQB&::(\ T@ 
@0>U$BH;IG;Y,>!#'*/'S(+''P73)GC*C&DVK:N7>7P, 
@ .P205YE0Q&9! ;L0%R&$V*"(OEG/LH$5/<_!3F_<@4 
@_ZHZZ+(N(8XTC*%6DD54>X=+D#)\N*Q^>6]>43T$ MH 
@_1%+6+9D8I*=ESD01S;\/9;RN0:_[X<WDG;:Z_,)<^P 
@*JA(*[Y%@8F%X_QH"0DE.=\ES2;_T@1(O>"^)O]#7/\ 
@W,KSN4]GAVZ9  &,?_DXR4^O>9J'DSTO-7S.29\T5F4 
@-NZ(#>NULSAL,F0?Q["(YU:7UQ8E%\X;LA\"PMH]*+X 
@1JVUC,?N8AO>8P"/'E(!='M'X,#K5@ 7&<RZG'&/]K( 
@JO/-/Z#UGUTAR9X0!] 4-! ]X$YHUIQ=6**62CWL 9T 
@#%+D/QR^,4(DUBKZF0NB33.$/(;#[7)U+,\46SMFW"4 
@V7]DQ1:$QY(AE@7)C.33Y$1*:OH;>ID"RYG^_,/-U_L 
@B=B8_*F@=PJ37"+"4K<[CY@,DP/U_S/6L?!.O#E?Z H 
@CA,.DI^0YNA?5N#.K,2'-&RYF418H2#+6"9ILAN]=UH 
@XK!!X ?TM8_5V 6IM0_&)>04'7;95?ITV/4P*IWZLO8 
@ +AA,ZW<0D4O#<14O^\9YH]45"W2'^"8;)X?O!%Y]9D 
@/K/RQ/&EW+N\P9I?SU,I#$[CO\J4L&@8;J _C>S$Z'< 
@+52WO"T26A.;T^"BD6 BEG4<5<F<L=KE4$0$*VX7UY4 
@%:0]27>0+=Z/)9H*6TPRRVVG_AA <S0!]Y@O[N#G^!X 
@$4.O$D 4-.][Z;\[(.&(S%VVL?8*X(H/*-*'&V6 "OL 
@[WS]G]-J3D-\V88W633(&<M"G[M*E4_,^)!5,9RCDOT 
@;"]1.\PIY95I -]I'4<GQU25:=<>.H^TH8JY[K<9ZC, 
@V]1%4Y+]KVP!'\H2Q$=<!GN,A U5,'UVMYH<62W.RYP 
@ W$&?/.U2/8EUNLBTZOV2E=<> G(W4F$1F5 OQS.-EH 
@''K<_,: $=,R%D26_S:2,N[%-,Q@Y!RY*/DKDU60<WD 
@XP&HJQ0-H'CODNO6.IML'U^%'Y)1/R+QN*7&:"T%NV\ 
@6 KV"F:]^0XM83\&CO69==A8>8Y7C+&,3U'^8&COITD 
@>VPS8R%]*L:" <(N1^ ?F7I1;10EIOPZO#,6MMP07X$ 
@ )G&,Y1I7;%PYXXK(=X;_!,< V6,<N?&TFS4D)= 1^@ 
@?LNIBMIH%?Q3V"(X'&G#]SQ/M5+/?,"V_MX&G'&Q),$ 
@]X)S>U3T9)WTQO=F)'6T#J-W2;>3@,-(X]FKYSJAJL4 
@Z" 2^[>F)\GM#+'9EV,"SF#K+9PR;P/AN@BIJRL"A!P 
@1AG] N+_ SQY:+>L%-H.PW65@7=FR%.:NW<NV^C1IA@ 
@:E2ER>$1SY$Y[B,2PID;%G*9C;/6I)]@?M$M8@0(P[4 
@HU* A8B_OGIP?G'3R0NXU]D'U3%>QYS-XX4-!O"RSW\ 
@'E+WRULU3X+KN-SI#P1^)G.D(&8ME[4/OQ,;7CNHHZ, 
@1J]79J=N<+*G*UYMW?<)(T8")XXE>(H_QQ9=G-Y!;'\ 
@18ZN+O9*0+12SUD*-\OH%MQ#3]<2QX3NY@^9"!J&#:$ 
@A!S^U7 +$&Z';,0!Y/COC6[R/^_?/@VM4V!G%.Y]'84 
@U7UTS_^Z\/E;4-:IGEX(T*C58$Z+WJ1ZYNXKMRB-=?X 
@&NT)0$59[L>ME+PD6XG)CGYCU?936'[F3 L]PZAG(:$ 
@7G$% N&^27]0$!* $<7)N<Y_^8YQK"?BHVF 5%^BG08 
@#VS7<7A$!OI6+CNAY@E*\BI6XOGYUFA*?%TCWLQ.U14 
@8["AK\!_5$P.=:_&R*YUN_@V%9(-I?U CV=ZVN&MQVT 
@MNN((?_(Z7)AQ#SVK7$@+KT7*LA#?\%O*!F!1L 5<=8 
@'8R(9*NW%$!LS$1^ 0T_NE,*7N"=KE'5@?/Q6H .,6, 
@O\HJT[:LM%&JTAT9_7@^+ZK_(N.\?#O>47A (A/T)"0 
@CP&0E9^(8;LE1!Q]\3E]_"JX5VD/3KH/JR<Q; 7YOT0 
@T#UJ&VB+(.-LGS#,*D$[Z1.SN8;N1K:\D?8J30KB^K4 
@QBW7:XL7C0QDWRW1)IK"Q'EJ<VD,>_1<+>&R!VN,[E$ 
@?*#M$^^S 4B5]76"'?$KO&>'I^F"<G=OQLN'.S+6F>( 
@P0C.<<381T,A6I"_"<*#;@[_S[*O8U12(- :1(1 2Y, 
@Z.3K0I1;Z@?[:)='I50^VV^-;A 3_8M7V.>#"&IKNPD 
@U8]\05IW)NZ(N*E_G6>)RS5+D;-^BB7@&M!@"7/P "\ 
@C'"@)^CG)K&':6!>?.Q$OGVOK_Y.Q@X? 22-YTGMW.L 
@*@L#?22):5:642[HQX) )2:D6S]6^PWJ-)@^,[K[81X 
@!/)<H6-*O?%JB *5_).VXU#VW\3>\SKM1G/#FYB.Z$P 
@N_VE%;KRIIU%7N_^%,$K*@!;<'[5=]K92%VYCM#43/L 
@M0TUD"7LX9:A"F6('>_$N2:?4["J2_N>-F#_R)OBZ'  
@442'1;>$Q6WE468 701]2:,VFPN#_(/TD @J[.=*Y)< 
0P3:V#4; 2$/P[J"U.Y4 7P  
0'=^5SJ[_);-* \Y-**Q"0@  
`pragma protect end_protected
