// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H_6Y07^>;5YLSY%;]8&USPGY1"QW$Z\D_<U;2N^VO>N*X-HB2=G779@  
HVTL-O) ]CB-DL4A!.31'\8)@U<;O'/-0*PJ$&9DQ)XS.U>>O2(%?$   
HQY,FQ_*E71K@"53]71E!4*)O3;K%2#<7^H,37GK:$%QL0CFQ68+H.@  
H8>NRMC*&C[,"'2>)7<C1\SQM DF2@7R.[QZ7H+3RK[<=*28$26GX;@  
HO>IUP<_G8&Q2:,W+&U+0B0X]RK_@@E<):YE]NIPW\_.3#_>@:96BNP  
`pragma protect encoding=(enctype="uuencode",bytes=17680       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@EK(*RN\U)PGON/H$0#+F^Y(FJ;!15@K!,Y:JB14KAQ@ 
@QYU33-3I^Q14<\M.'LV_S4H4D(AG%9)@HA'. ##Y'DP 
@U:\W9UKGW0X7O)XO>D%)!A6JXN0B9>4Y@/SV2-\C%%T 
@[,#._:Z.]Y'^R:#ZU=<V,H8AC)]1>5,#*:)<523^ =, 
@GP!^X>E\#"#-9,4QTJE%<@XZX>G);3!33@[N%.!O$>  
@):SVBAL*KD'WY>ST_B"5Z :FL,LR3$,.=HXSK[X*Q.T 
@^=*YK"P9ID1GR0+,T$II1IJ']^M,QI5(E,:+8W=.94, 
@HT\>U>B?]AN:7Z._%7GFO53=1:>,ETK4M3#2!XI^.:$ 
@H;-].@6IX''9X3@JZMX^KI*0?R?L8=H"R ?&_A4E)+< 
@^R1AGO5=<9*622F=].D[:WA'_2J$;<_)ZC+QH>X2+JX 
@IYH [6!NR2!$G63H]5;5*T=[/:25YGOGW>@-%[,N<^4 
@0^=U>\N2;Y#[R%!PS^/18Z9C,X$!$(4DGM@YQD+>:20 
@7 DOZ4*HHLYIR-W?0@\4([*EU/MP.2Q]'2!^I,=<*UP 
@07WXAZ/8,8ULVW4N GCN<?R=K5&SD%P8.J]E;-@% C0 
@1-?&TUZ)V@4H/#9"F:?&5J%2Q"D NRF>BJ?9V?6_SJP 
@(;=:D6HWKB,MQHO==].!%>;46A=3CL#1U.]P_E\Y^M< 
@X&(3X1OL'[D5(KT>Q!2ROV%A+\E"$EBVI_M*G]X\N$, 
@&"C+65HX10W@0),ZD6HM%%L,S57XH".%,?T$_-E\*78 
@8%) F,.>;.^R/K.=!(KBS*ZOBBSVY:,>OL?NXP@IB5$ 
@C3((_$QX.:7!!H0*2%PYN)SK\=Y%\G'",D*P5S_Z31@ 
@ O_4?T!'I,7A?4%G86X]U(I-=N"#Z95A>XQ7HWGU;I0 
@V>8<;M'!0C:-=T/- &*@S)MECH]9 :YAV^0.#&/B.Q< 
@WA)6($8:D 1#@;%#5R<;W_JMU>6,.&%.%3^<+?&RO6T 
@\#N=W#C]?P1)V63^2JR.,'^(%S=(J38;,MU=6G/3.I$ 
@L82S/!UR,7FWEE\.?C< L^[*Z!*5$,3:2IWEQF%D<X0 
@T@3[KO'VH(R%(3GDVHY/[([77C\D8%BO+!;^DG(B!08 
@+"$ACK4M^V^[/OBT!*R6.RRU'"K2,_RV$E FM=\>=?D 
@(VYVIHW91.>8J.&UL+.F1GN'3V^'3L4U4Q<XG)UI730 
@2(' -TRK>K<&V?+Z.=OM W,D$ /]'^%@=M^QEIV_-8T 
@U217V@+ .I85OK# \N-^<B]K2M!S'-&ES:8NWL9"SL8 
@MEVP6SZ"=2]-$F ?C,;HN&*$Y%2C)_[4=Q$Z ?)TW[< 
@>BYDLI;I]B,0AT?$=TIJ[<QTY%FLB&<G;P&>>X/$7_( 
@1B9[EGR1)![03KAY)MF ]A*YF$M#(3W(DE%UFH.AB$H 
@"E.0 J-((?+HA8J*\R76@8IN@^9>^TTZ-0 "),E/'W4 
@H*&0#;T 1RO'G*#:"LLQ$06%]K;T_G$&A'_;;"9D*/P 
@2/_<RDJ21I)=&H(2@,,KXAY&\8Z]>8KB3#--!/,C6Z  
@9G_7.SD%;#2!JPSN.]MH A9A#F]D$=4S.JX6-1*4^$4 
@_Z7U#_^S^W_S5D8R.V-WA(.8DG7"0ZA^&9X:(6R;TV  
@,98@9013$@?RY-R_B3\N>;8V?%Q-*?(\\TB;2:O+WG0 
@]4LP;%/;"/$-.-R3/?2"$!^GEU6-DOY=D;^!GC=X3,8 
@0=\[-"RER2)/J5)Z4Y[-]AW(D[[:>?CK\A8>&.1WWP, 
@G)EJ@J+BE^U'!\U//6"Y?!76>;%/Y?!IS8N2>T'NB6P 
@0>Y!,5^.*IPJEEHM;^I;II!;3A;U<TAY<;G?)L7*V_T 
@K%-P"0IN,GT%F6Z8^(1K\'SA4"YS#YCO?\!)&9-^!;P 
@JM4CT]%.ET)&HJ%/HC$#[CUIA:L?N?M^1'F-,3XK?!@ 
@'0G:M=Y]TJ;!AQ4-<&(DQ"*/RYS1+L2GZH?&_O\1*E4 
@AX2GS;EK.XO#E4R3=5<SZI=<VMB98!_8^(<^(AW#&3@ 
@L:VX3$)SS68B\.?2KADZ76_*56A)Y#PF&6D?C^2X4Y  
@Q<)PPK4RBYE>8PQ+U#*T><D_'BS8:9^O3I/:#HHEG3< 
@VY 3 4G^D]<WWGSTL*RB)4GYLWK4]<Q!Y!&-T)LCGFT 
@]F8KK)\ZNI@Z[A6D-V0&LX"$/'<9IO"9["![#8GOCUH 
@[ET5\JP%E:CN[ CC>9:+QE:9>YO 0Z=L9W;'&%,5!,\ 
@?L]@[IXJ4'T0:;@'QHV.$]#=LR6C9?NJE9+FZ]V\1LL 
@OO+74/[56NGG$W''<0': 8*94MO?PKFN*D1?_T3R+,L 
@ %KTM&=)9>*^8R51BQXC3]>FLJGBM>F*45)L%=D-C%H 
@:&"TMBXRE?Z;,L[9-M+2N]6;_-S>A\G+_>_,=22M1%H 
@.75PBO9F1P[\\R?".)DMFK"?A*HSS1A%",+_9C7%'!4 
@J^NC35M-0_Z2/3B0\48 9Z-JP6K9]"U$5.:959/R134 
@0D3:+E7?!P(!V1]A6I-50JNAOC<LV7JVYZ?;TN^_W?8 
@Z/[DGM,N1F4C9X3=;;IB@(7!F 9<W1X[1,0=RIXU.F\ 
@8-=WJ]%TWU?>&0! 6T'#"O%3PX:WR:W_@[KL5^;:(=H 
@CS8?HQNRX,_85>RG<MU;]]J?![]0?J%!&XF;<>#NM!  
@:7S\TEAT%\%==JUREUHL:,F;_[=?X&.W G5SGI:_?)P 
@O/S1Q22NV)Z4%W"^ Y>8RN?#G6%K"P^HZ&)%;>\%S(( 
@1&^)/=  @@.W_=^+GGWI+4>:T?:$RIVOCH'/H-CZ3CX 
@!/I._Y>$JSH]R)0$\#,:A*JC5(7O9*86K9K"M"5U;.$ 
@ZB#A8Y>TG%Q3!?X:1I%RB"@F[KS,JT871D2C8G;UID@ 
@#FJ]_E77:^HJ']51H #_M-@U8?\/JR/?MDX$A)8OS>8 
@HB2111&1&]RKZD?-7S@D\-GT -V*QG.YBHDD,?2.,'P 
@U[F>+69)/UR-NG/@B5A[J#UCOZFO:?B=:$<U'UK2KK8 
@,4?EZ 7FGY3>?S]Q!WP65/KA^00:%REJR-"+K4OZH@0 
@'-LPLG/@4;KR[,?N1.FA,Z?SV<\+X";K3!5M@&6NRG0 
@I!.EM@/4>VWIGRX"*J?[K E.S\S*)YJW%0*6XIZJZ;, 
@T6P'0!5  3<[)!E3-$Y+-W:M=QYO6//(4'XA1TAH2)P 
@S__&!4&6S#GY_QY)#NF&?S^+=XJH+Y1S 0?GCP]=1'$ 
@DESPQP^0??=MECD-&]?G60I@R;TG@*A+,K2X%5ZT2B$ 
@?2PYRX:7WT(5=IU+COQ-XL:\(T,$\AN>73SNV-6<#(, 
@R+9U/!0)%%ZBLE%E(^GUP?N7WZV_FM,"LHU>4^5Z^%L 
@+N;<((7"WK^[[F)07DI^E*ANYH]>!FGWH&]'A[@AE6P 
@BX0,I1O7*9K9SIUEZJ4:1=M1.JJ-FF>U%S_ _Y$I)H  
@G D0=,+TI=3?*<L$O[-XZZ$?%[_,O?;_!^9:=;_\3PX 
@0BV$"%E<]EWW-I\SKQ[2;H/EAY[8AB-/M!J''CW/+M  
@X[<,+)Y\)DG9USR27#Z5?_WI:C\_IT1R]QE?_/S6ZSD 
@>4EZ9]O<R3#?$ RL%>E%+-=TZU3IX*H'J&TX#$)_Y#  
@3"[S:I4;0TN)FMP2A3N+/#W0)9(MMB6BA"4I*QP7T H 
@6KX+WK2'[P\^==6D*)K\@")+[Q867NB0K6TB"5-D1-D 
@H/IN>9]>Y0R&W'SHOI+]:0:.%499B=$#L_MGC:"[8>, 
@WEJ:?!X723])^&S6E:M?,0B@U2!'_;JY++^;4HP6W@H 
@-)J(98*X%RJ9/41+P7Z:2>F<,;WQ[*& %2BV:$II>2D 
@&SR%-$!+C?./G*]',8$#51:MDF6#S/GF<&(V_C#;BL< 
@E]'+$!1FT^4-S5K&@JXJKN2IBP7 ;70H@A13@/Z_V68 
@F 5B;JM_8@LEJ6/ %B#9[YZP5K/<2?0-WK,^63$D*Q\ 
@R^S3B-@O<-N;*FA^T?71^=;QO "W+28^PKM?0*$9.<$ 
@E%=>!XU,>GUO .M@(3>+^"DY_TS@%G]"35@=\3ETD]4 
@B*2E#TJ*4&UW9! :#KPE!/WF=ZBH'*B=N< -N.51OQ$ 
@FV0PINH;H>-V4>P-$]$ 5Y+?#B<;XJ9C-4#ZU.)#\!@ 
@6!$OB:I2V[(:/$.DBU8^3>RG;G$KR-,GT](OHQO(U+, 
@R(LV!; ;:LSWN1S7&V]=1*@AJ*BLBZ4S;U-*,A_HS=8 
@R-)H+;VH>]$T(6[$_N>  W8+0SFI9A+/Q1DTW$'@=0T 
@#]5STI9[#%+)F0EUZ'J]3P90\*+_I6-V#H!\EX%_Y.( 
@^YM_I[5/U%PU)D[<U@%I^0:7@)#,4=,6+.%)0;_$9S< 
@2DZ0$IS/X**'L3IG8-F7ULFSSN5[0D"LE.K4#'(K[=< 
@;6"<F/Q73<"+<YJKZ;\")'45(Y1;>58U_<\()[OU78  
@81$=O3>BOKGHG H[I\HQ0-N1^N%VH8'5**0JK!#?YCT 
@2$M4Y9:X&6 3MX/7A?I(-V%!01KE0+'@N./5*_;RY[( 
@:0IYR21@B-1,R\&,:>%(<;Z2TMRK5#TM[]XK3\$&L6H 
@*PX@,]^?P%3J9=D:6,V6[3<\W&!>@T&_:*^F7=+ -7( 
@*U^/1?\_&CZ@%F:*VK3K48N8J67<Y05O,:#DTHPN[<@ 
@7K!C0,2,#"-6Y0D6;J6^)+_"T>-#E'"[3FSG,C7UP2T 
@\A$RFY9_$+CB0M57U23[Y>?AOO3P+.$^Z&&H>*_;J#8 
@N^X"-@V"9B^M!$@&03IF]+?K;SPU58):O^6\8(@>'CD 
@IR?R$&B9U37D&T=("<A)L8M_[T_3RL MF\)]3,I"&SL 
@11=+A]"]/SM')U7 "072>MUR@WY%/#^H[5WZO>;1GA  
@07 4>Y9\F-J#H;[?!<1"69DC0L!4;P/S31A\J&2+#,D 
@QA4J;VH_B+K]"K"/_0Q!WB%8,*71?,F?&QR&NX>MA#P 
@@Z&1O?J)IBPUC@(!-<RI;>K5FHYLHXM@G=*!':DXX $ 
@X"\$@_JD=>@@F-L<\'2ACG491V)?*?/28UDNW%&V2   
@3EH.G#O(EW8Q0.#A#>C;*WO@!RFVT$Y^* +-;78D.#8 
@G,FS\*L'4'M^N774ZZICW[3EDF%5;L@A5:ZR?Y.-P"  
@R3\&?<;?%^A>/O1V1VEY$'T&U:8O5;AFP24]D$P2[EX 
@1K*.LG&RV:$B=*A653$*0G:N+2QN]<50W3<1@R7=8"4 
@1;9$0_J:4O)O_[6OI%4LU <:0+)(TY(^!'&BR/H_;E0 
@.)!%FNG*Y$)+CCG>?U8(K"W42#"9CPZT)#2?&2S2'HH 
@G<;@#O9E-U8W#A3XCN AB9,MN"QU=UBRNVG"Y_EY,/\ 
@_ B3H, @BL&HQDI6ZU:AW$^F@E/^<_WXU'$T)@<.A2H 
@5JK-N)4](\V9Y_%X@DE(?C,;]F[22/G'X5O<!SSFQ>@ 
@8$OX?Q8K85RESCR[T_G8CE?+,@2=C7/G+\97" GR4(4 
@#=$U#_)\?;NBF1I%)>^+WMAHY\ 8$S<G$CW":>S'!>\ 
@,\V'<V3O";'WJ+#Z>)*A$>0V)2=UYQR$_ 5M<]SSL10 
@US[CKO,,%!]DG@!*V^;3:+^=AL4H;[(V;YT/R[, P,P 
@7'\/<N#P9ST&)[3]GYL.FCDCWR=W%(?X5WB],6F^]M8 
@,*324D$8: 3=@S/\RST7H&M]JUQ06"X3I"%,Z6+F!'T 
@/"M-FOEE2 B4$'2Y>(P4Z9G=3;X/SM9--!R4M&<VQ\  
@UI'2KQ+K30A<W<,VB[4HSW;F+ABGP2HIXS3*F97H&N@ 
@1V18<9,, IL2G7RO&""K JC$1E %RB&'>]&_'0T_B[@ 
@!*' N!SS%Z^SNTF/ZN@E(]/-B!P!2F /*0ZA;FBUZ%8 
@P[ T"X<"TT*[5=-TY>EUXUELM6S"='LS#RYSI]<5;N4 
@KJEI7.0A[G0O@5Z"/WX7.;#%T?GF6\XWXDR9#2E$R0  
@N"D4&5(]\FZ5E1@@\!@HJT=@4QVE%"9![TU_@1<3TBP 
@QF @XSEQB!P$J%QQGL]\6$^NV@10AWV?.Q]S0.KWB9H 
@*]@\4].]HZ7#6F9UWNPLYC=X531> \K\OP7_]%1''"@ 
@FX$W,/XE$5%R*"^@J['6"7+R=I8RCG#:JOVTI_(4"]8 
@%8[@CO-2SN!,E^8'&\C5GT#H4"<3-DOEI(@/19$#+QL 
@]G:>.ZXT';V:CQ[0BVE($1NXLH5#:!>4XN/V\TO5LJ4 
@A%P8[R5N.JCN\&D^?$>%MZ,IA0G18?W=A)%>TUB;&7$ 
@45RYX(4POKJH!2$&?W! /4&7X#OD6I=71:[%".0]ZP\ 
@1(=57A2HUH%#BI#;QZ$6TGO>[U>;AM/\#D_"?:Q)%Z( 
@'K*(G,01) <D&K9S?0MH\NL:X\4M2C]^V"M=HA<D)>X 
@1\F?+49CYBD1%UK 5=\#+0&^Y?X6B[5;F'57K!H(>'4 
@3=6&RZ=B/5+72>27XAXD))Q[1/K@J2$0'FW]6E9DG'D 
@O()7>*[F]3()\7SG ?6.I]@8K:>!WC?;(,+BOTE)K20 
@"8R2T+:8JH31""H/,H$5M_PG8!\]#'!-)M'M;0C [%\ 
@.)!8P,14W5B]VL'[O.U0CFM._28VA!*Y\MWD]-QT (D 
@$*_('ZC^=ESF"@&I>?>D@9)T5P.:3+443G$&"V0AQM8 
@M$3KXL8WK%^=("@SKZ:R0DB?$U839[\T"A7; M&$R[< 
@+RD&7\/GD'4LJRDV$;TE1,_D;>>^^!L'R"-SQ@=(<ZH 
@:,'^$6?!I[_,HNK5)Z8CC!O8#L ]VL437#9AHF,FS?P 
@6@A=;<Y\V._:Z7MD$OB0[P/\,;I-I7"=X<,&T'2HWTD 
@$(1V+NFK7X\]\H[@"1-L-H55>08.+X3'RLL<MKB6,2H 
@503[%HH2J:]:O11'@1,J5=3T4?EUX)%^GPKM;P>;N\  
@8C[ MXE2C[8G@8I2FPC*=:N]=RDKC[<$/P\<GO#SUT  
@!N6+>*N1!.T+FF05I)BR'I]> ,5OQ&:/=#"VYU(A;5@ 
@^"^33]>8";0+?S^H(G[YOT5Z9D9U:GNEV HS2WZ!5Y4 
@:[55NJ57(*MAZ2CM?M,[.N<R*OPG;13EA;Y2OG'VELH 
@TYH,*@3ITB3#A"=3T95-S%]P1T)#3!ZV-&M.BEX%194 
@DG>B'6-RVQ'.2_]JM.\K4CKQ( F9Z3U.XE=K0./0(+< 
@J^4^FMJYD6N'[0"JTXY('B\DP3%];PF@(-\YA3FW7OL 
@Z_IEOW5Q*Y#7'%H/>6X)68&,35'MTY]+IB8PU_*RP#D 
@YNR/K7E_UW/Q%7DN 1$P!)%>K3B%1?8\WLJW64>ZA:\ 
@B"*'<9^'#]V>QR40Y%RDEI#]2SX"TTI,^L4T=I^\'Q4 
@ B8"G_RN$$T?OD[%#73F)472&F  CA:D#7O8L46R] L 
@EK/!QM?#^GBV$2'UO\K6],E_V6Q?+7FX3.YW(!!O$U4 
@S9FN+EA!/G[DHSK>G3D0E,.]0277OV"F[I&:&5,B(?X 
@D9Q910.\V"//5J=G[0RJE; [-#ZZ8M-9S_ U/U [O#X 
@J_>]U%]2ITR*B0#0-4\FR$H*N^7+-DX%AT-_"!6;+7$ 
@DM*O1<X[:M16,DUYB\!/XF@OA@,3["0]^.395U_*%#< 
@&,O>IWR23I:L;8T^>H@O#(?GVFL\\9;-IH+,S+V%1&0 
@W.2.&+S]@-II@H0_6YU3@K,GV%S3 9'JP5V5G ,#BMD 
@#;3)*-> !_@0,A.52)Z!Y.WT^<X-:$1__A1[!^33Q[D 
@K !,&@!>RL'Y>M8U\4$!ESHB=FS#/N=&;&!S66&5];\ 
@%%L-@ 6N<PZ&6#$=WZ5A?T8MHBENF90K-6FW6C1\$!4 
@(J$ZX@J,%>OIH^&W>Q*[@HCCTWC[_I@8L]!CP "*XR8 
@'KH"D@IH&% $(Q=R.+>>/Z!F96U+!$<'6Q)+=.L7R+8 
@7E2M-51CD5 XT_P]?DBN]%M34LV^!3WIDO()D@V=HLP 
@MS9)>9MCE,^PAX2$,@@DG4J:Q@UX]T.YV"]M,=KO$1, 
@!8CZ$,^5MZO_#:S5:+ *JN2L?F!.L9L=<;$7.\(RLJ( 
@57*0U70]F6.N8*;^4.*&U/&:C>0+'^C6>I0!G2<J#%X 
@'H!_FV1+\2!)-7R>92>RG1,2B@G5,D7OEU#R,P\<L_0 
@Y(O I?JTJW5"\4@0EX-:NCS536I.%V5(\/PC0J#"@(T 
@(53UWH+DN?<,FFG6=1EKA&ED:(J,K*&;#*$8[8Y*O2X 
@&X! (Y?Z^6DTQ4%SJNLPRJOP;"I.E"W[U/_$:$J;_UT 
@VCO,O<WT;X@D=Y"&!2 9@CK;E9FAM8@E'>[G$<R$4:L 
@>,/MAY+Y<AC9JT]4._0"X@] VH;Q&7O![V&%=>Y&A:( 
@&9X[_FP>S#7)A.(&:5*#7I&SD<LMN/(.=QM&R[B:F0P 
@*6R;S9(SHY7-L]:<K?RMX-ZK*^)Q:@)H@(54R/RPE)$ 
@/K4S:8IIV]IKYQ*S3G&[D2']\MIU=9.RQTXI\Q=]C$4 
@]_R!7;+P!SXQ%A7X?WU4Z+8[8@"EGZ(GD$D?TW&7[5H 
@AG2*BU<%KQXG-F"4W[(Y>=2DAR5W*/9^$\UDFQIBJ&D 
@/^6TX=#BMD<%P_:,WF,)Y21!Q"\23?'>=G>M7GIH&A8 
@@<&]Q5*1ONJF5+#M'2[SKO.MECZV+1)(G@VVV09,_]H 
@K*>#L.K\7ZI##"K%.E9U?,0YO(D+\;/-SK'M)<(D:0$ 
@KJM[*% :9-KR#1GI>D?PXD!H/XVP=>B??F\X5MZLI(X 
@3G@B#0)DUWU\V?Q^ &.Z,DFQ)D-/ND@H(!G*=TQ>>^8 
@C,!,$W [R64B97J+I/_=G)^^*%1*4PC\&5R'0<^]KQ, 
@(9>7#^OSK$?ND3]=('6. $BT'9YDKB';-IC0+'3-^WX 
@ZK'8G(6V%V*YQ%])8V/\> -%$[CRRZOOF>R>M!KHA^X 
@U=&%-'YUJ4M^8R2%K*12IW746)O"!9$%'^U[ZZ/C4)H 
@.S5PEMT8%PG.P_H?E0]L8*E6S%1NZ<%TVH.TT'G,4%T 
@; EQ\;1"F&QAY@4:/QD:EQ%]M>Q4_(($0B&P2%B!X6@ 
@VY#9@F5H![0Q2JEC2 J?K$S\" [@J+Z?/"%Y]TF8+5L 
@>5";,J:S-EE37<'MG4:/P@D01'P7P:Q/O=;,%T3=**D 
@J[UL*@[GLC7*6@M5\;?TO_[!]>"8>@MF:RGCH="*?^@ 
@K:]\^F)HTZO:2?X5YPM)8*[',1-3=W]$L.AOWZU-5>0 
@J5VNA31([[9A XVY)^L]3WD#G5.R XV^DJ7KG=(T73, 
@,C:MO9+[*MO,ZJKU*MQ^%C1*P;RD#'O#$R,"(@FC.TH 
@YF1QAC&@YK(BU=T9'+=4$_^B)E=M&^UWG/T ^=_AOVH 
@T;[K*PG >O-7F9\'Q"5)ZKDX0#TFY WO]%=4KQ-LTG< 
@&N@P""3!!?=9@JG,[5F1^4@SZL+LW@S30U-D"\6VHND 
@+X..M"%.)%R'JVSMJH&^1""C6P*[//*W2TL>H5X;_7$ 
@OS:RMX;R1_[*/A\;_"\KSUQBDH(%60%>(EL(T\!8[Y@ 
@&!D3OG7A0&9;U \F<U.D-]C:<&MQJRMC1WL:$96@:<@ 
@5#VMB/DO@*\<&+A)Y%C*Q."2-<6\<$UE%LVO%B9,L9, 
@$YXT2R-(FO-FQW/+(-6IU6@Q>Q;SN'6KN\S#C#,+)40 
@).I'YC\W67&.>C]UQ.D[CI+'SLS7'@2OB[@V4]1&.%  
@4&; X!Z.I!2#',]&RSJ,%Q7$U0INW*PA3]5X+M8 W-D 
@;@+C(?LF"E,\-V=1$+OH?$%9H5#$D:6B2F-K[;R:W$H 
@!;:%)V)"Y.K%W#O36*3E.R# '-V\&1M"=PVE^D1'DGL 
@PP%.TV6,(3/&X=9F.G6#KU;4\M33FK^"E6T-W/\0KHH 
@W/$2"K]033WE?:B,.EKD;72H)2<EDOS@\8CL577RD_0 
@-4M%@ZWV-_[;M%IM>,^3&A'),L2?6'=@B_-#>62"OJX 
@?(5ZX&ZBV\L1M^_9(ZXO@4U!E_N[WX+4G=,%*X:[IID 
@88>"QRQ=6>Z]OUGQ]6Y8Y+_-4S:?V!X4<NG,; Z:Y*8 
@9W&AGOZ31.HOIWX+<3/ VH__>NCR\)W2LJK!R_>9+.  
@SOTWQR.Y:%C82Q==!\ZC<H4+O@[HI3N<T6M*]K-Y!28 
@!IGZ!!2$\&4# _=FV'R%W,GB8M-S'L+-7"L^C,^#IZP 
@,U3;#D[R%< [<]N=2]FCH/T$:DU_-(G&NC6OR(PC4,L 
@PQ?1K/O%A_&FS&[M.\(#MM^/JU_ E=/T4 .@=D8EZ)\ 
@@O/_+*)DW[9+?Z9:D):4H+3E3R71"@6)D*$H-T_L_O0 
@+S#>K5#PWP+(3F!H"R;F/7IG7/E+J6FU=SXUR>!!V9H 
@Y+B=COQ^1C.%%E-*7+H^8CO>1.Y2)0#C9!EK+SU*8,@ 
@V:_ )\^X0;NY0Z]9']J8%QP]>W $E=#[-PS6#3J64/< 
@J1)W"L5_&P%T/^WF]1>=\Q2U"ARQ:\A"1G\LZ33J&4H 
@S2,9K48$\<XYIP0<-CB/2'9_(%].5)=KXO[BL)/XZK@ 
@"YC)E\J;_73N(67[= $C0\AS5_"[E8;.R4'M+Z/[5$< 
@)W #XU91#F# -WKH_4UBZ?]+N=S#%]*2S.GH]EW'KG( 
@B56Y/KL;,9.QT4:HW]/ HD5W9QSJNB767:[@WR_P?]< 
@*.+TB=99HS6@@4T#>^N<FFZ(!]P!0MHV#!"-'[8NIS, 
@?SMZMQ.#89P^'-5\[O<7%EP#G[SF<U'UWO@E4[ZVS<( 
@H\8+%=E[_89+JP:D);_MDA3Z#G>X=72Z$V^6ZT'.UCX 
@/[[I>%:8TU3 K8),O.PI<;AU .D?1,U)#MF&GW!Q;X@ 
@-IF";/Z=>YC*#,DY\G#&37KLS_/[?6G;YWB39V>CO]P 
@-\*!#8+@[-H01Z/_8$3.BX&S!8 X.U72LP^JT]/P3.D 
@^1[.K<:]T*I$V>&%SU0_#+3.V#>,)=*IVH@H +A\.$4 
@P'"]]O)MH<Q'QB"G>J0AIKL-4: :M;_7]OPV'Q.%=6@ 
@3B]+%F3NI6.*+^@(#LFZT]#F1K?U]K^$3F92'(9!-A  
@AI]+F Z+)8[=!,\!L2SHA,/_9OM:,'J6^Y++!EWUHR8 
@>5_.@[U]K3=C:!7SAJ"0;)4A<N^3^O/+:XDTHAL;T+T 
@K*#!0)>V(C4R'IH8W%<*SR\;=:C;O_5;%W=3])021F( 
@XWJGJN:."=;V4VD:IY-ZXNWH8MHQ'=6083S4-)L=: ( 
@OTK+Q;-JD97:J5->9Y/BO)EEE.OR*=OI%'I&P^(,>!4 
@P)L%'IO[JX]S,VN6M9T@7(UHNY.T."M,^#B*[+[7 )\ 
@^P]<W?>"AR7_(W4R)PNC[SJ8Z D6JV! *&O[#<KK((< 
@]4NR7 U%]PY*J<+)K # ]69/X3$=1YJR$0ULF2)\91D 
@0\OH@=)HI9*NM5;3XZ/7B[N^>^E%XQ+=AID"V(TFZ-@ 
@5K:^0W%)AH@]_85!307;)D8?_W_9;IL6=J824F7V2#X 
@"$)_\.D3!\BL4&AN9'736@2JAA21-.)FBVN\-]VCUM8 
@V%+L\.<)-*RH:_[?%FFS?(:$^(4\4GQX;.F\=\&NLL@ 
@X0E:0="L(MBED!)1=K6R?0_B(6 J&,L+T!3*O\%%BD  
@=,W,*;B&""SY=OOKBFBWEF"2Q4&1,Z1:$K",TF^T!%8 
@U?4#J'U8V/W%%)VM8/J;.<%)U&Z?F)CP7%S+[;%V\*T 
@*+AL'^$Z6.<<KB&@$UGY4^+1KFQ!PL37P*CY39P^T($ 
@M8<?M[J(Y6M(6KY)#P0S9@Z*B 2<C?25@,[7&K,*>&4 
@9>UY61V#9^T&E,8"T2_&HH!J[, :A<-O3<5R$P3HOF4 
@Z7JYOWMKQE@$^+L#<L ]O0FVDK.$<<"I@.$/-?#5B+T 
@J/^_B,VXQ2<R=!_7$S7Q+H_HL!,J).121]&@O?O?%Y4 
@AHA(DPX-;S!(T!".FMA]A*^8='K0#YW&E/#?YC?6M^X 
@+UJ=K:OIDK8<6QW\"/9 TMOD@-&J_,!H'.X4\;E:4[\ 
@:E_G=^,/F#5$\/;E+<%^6+J1X&EQ0<M9^\WOT F<_RP 
@-$IGYIDP%I2>9F78:WA<"N!T:*-%"O4B5AD5$F#%/;, 
@/8X*7&*G'!S$$EHSNU(6[O$M#%4V<E/,,<*4*M*C_D  
@.T51;=%%W@@>D,B"^"\)XD78X@[FK^^N!D/HR--$+W$ 
@KE;F2B-OBDITO_9"Q5;.(]C(B5YKA']D<UG$K%LQ-*\ 
@=MW:WZVNC6W]GO&*;(D:>-)F-R%IG&U=KJA<4!1"_6D 
@ \$T?V@@.U<1:8ME(50=/PZ\3,*IB\]6?:'\T!:ITO\ 
@" <L4_RP6,!;DF8.#76$_=VQYCL?EP&N<<Q+B1_>E$8 
@G$.6: &$_2SJ^\=1[RI.]TY*6R6('8FJ[I)ZL0O8NV\ 
@C3PSYF#H+FY8LN4*810DWG)_6;3X^ L5%Y*W=[ ZF^0 
@54$][&!+#3@T,O* BC'DZA_98T[I?'BVR5'Z+97/'-  
@=M\7"&A&]LLL!YHE&G)%&<1"^P9G&>_:!58*3+("Q@, 
@$2"O[5K^$#^S6LE2G;"A4\,JF\]B0OK= 6\O/? P.6D 
@N9^AR[\Q7L-D,+V=$-_H-XC>SOZUK0DU48XIA'=_..( 
@RY'B[QU/VHDJ@A+K5)N;T-6$W-*B265$W/=WN0F8,M  
@'QU^1%&,4BXH2=:]OF'WD9E):EM>3+@R>E=GE<3YMGP 
@KI!2)Y!A*%A T<RIS_ PO$"%-;K_9'WX6BEK[;9"_.@ 
@WD@:T]IZ9(@8*Y01#?4*+Q0T9>Y,#J8MI!_E'QT@_'$ 
@,K?; \:WWD3:M >>0E"',YZD0VFI_S%<58E-EHB#Y 0 
@*QQ_V[B&@ 6X-GKKA^Z=O>GVUD)7AJ(T9N2*NZ;^984 
@7^#=G=B!PL0))01"/,5@(SS9X<@KRN"'Z<*:,[BO#BD 
@!*216NTJL&/:  H0(9N9_&5)R/#<;2N1/N\P\ E##G\ 
@>EIM2T*@.J0XBF44&);23PWJJ^YX/"U>W_<-6=\X90< 
@!3],PB+I"8:"XQS$ 2A-]M'Z37BTC'SF*'[.ILJB]K$ 
@\CCTW<67>\:EF(0"N]5YT>N2E<9-L) <ZZ31]>HIXLH 
@&<NA;FP:YZ%UP6NF$C;[0N!^I+;V0TF09(66O@!33U4 
@0)G (TV3"+1#&M4^!A850['7PSK33JH\G:NNC+059<H 
@RE>@,.;:W]6 #)?F\7Y;($CZKFJ:NTCJA,OK;;#*V:\ 
@?(#_U#N*183N;RB=Y6=$.DK:EBCKQI$Y<G\D3.C6P1$ 
@V1A%- +]<IAN#]2\=('O3=9>D%2T&C=SE'@RO+T<0?P 
@G$*ZPUUE<J3EUOR*D<4=[_D?PI!VW!),X9-=_^_AUA8 
@N(L_=PKA2,;/\5^M_<G[,TR4KU*2DN>24LE5OS&:Y/\ 
@BYH 5V.PLYD86+'$4^:]C.!)0T6.&FFD_H8KO3L%7@P 
@*0-D "<G;ZW>[!8A?>B6EK3HV2T8H, S #;CS%WJUB8 
@[.&G31,*>^S*X<H)7<X*+#;QR'IZQNIL1PKXO-0YLV, 
@@,TJCY7$7+? (CA6R#?.4,<@=ID[2 QHQC5S14/V 28 
@<G$?=,EQ7PDAW2ZD8NNSWU(3#IDLLGQDUT7$YQ2@1(4 
@?1.IL\K\W]BU")Y?CO$*!&EV5:M-R#/,X#?N[1.@4,< 
@[89M"[5+]?HYZ\AM;P"_)\ZZC$.IYPM&)O:1@&\#QW4 
@.L(:\C+EK*TJ_(#04:"0\<]W/UJ*ERZ\=0F2_DWEL;X 
@HPQ%&/A9MI:PLG?F+U,]\I->@4>^O,;^;TJ2"D O6Y@ 
@ZWDEH,Y @N5=X=IA- >2=@?NQD\=#-5S&#]+15#I:\H 
@\G+_@X*DR5K-TM5*%$W2YT!+AZP0EATZ'*O]EZGFQ<\ 
@#=[K1INQ0J8O.\ F<?Y$53/(#!.^L4AM@U*NO_)5)<\ 
@$MAO$%SCY7;_U?C)'19P(ON&[/*Z;)*&0S";XYQ4F@P 
@2=Q@.<?L!<I]?1V".3Q GN3H9R_E%P^NC1D4#S/SMP  
@XX850['L#!\;?[H(,&[PP4,O?A90*]AC:^[-CQ#'##T 
@2VA=.?JBH]7=555DP+U6P-7X+^7@*"I\Y()-82".*D\ 
@QF!,>)LBQJ.023O*9FB6?H *FIQN<Z,XE<N62B(%1U$ 
@J57X/U)2X?2;[=+7$_,3\21%=GYT8M"-]Y'3A=:7:(@ 
@97*-_7=6=IP&"CWX(WU#-CP#^F+8+0 L%E><X[>;0/, 
@H'S)QNE%7(J"-U0,2B6/&Q^E]<*U1#(K/B'VHX*8>T, 
@-JTU1;"W5NJ@$:H=MUZ3;B[M%D$ L8,C$DI00@3X"H4 
@8^-3R.H^PQ$FMDYKPV&"NQ$<&<+N3*;.064]+VSK)_L 
@-:_@?-GOZO6G*!#["3D)0UB$"L%M<&-VT::M%777Q*X 
@4$S[/L1TKZL2%A4V:'5Z&9GD JUY%T?]T<,XE_60"CH 
@9:,?SIG%TAA_H8ZDN(ZMC7&.BT2DW%VU273E.V?(?\\ 
@2P: *+48Z]+54$:7"U^']X9676(7VRM/^#QS%@JDG[( 
@4#A^C8*G3UIY/ R-/4?2O0Q@=RNIL20&7U6K'8(+,/$ 
@,MT2NF5)8W"%>WEH\HM7.(@H9H^:(?FMOI!% W&I#^X 
@57,@W754[Q/H3%.69"^<W<7Q3"\[D#( 8A='2$?]C$< 
@ROZRM0#WXZ :[ UBTPB3_Y&X#P=;^'S,_I*4NZO:<84 
@R8TFN#=M^X]]:7)/_5-? AKJ-2S'RJNQ])UN];V.E,$ 
@B_\#SW=6 ']RLN"E++Q T4GSD1VQV*O$#KFWKGO78'8 
@XV0V9*TIE:@Y_X]D='$"RCCSD4(ZL0'OC.7,LW?%8O( 
@>C*@<(WJU.LSV"8>D"3!=:$5*+M]9N "RQ8; ;P/?0@ 
@Q'.=27)%% ST7&)Z#%X3S7ADF4^%GX?SBD-3OH>4U>X 
@;B@**I*&%; R4*:"CCR",<0M"H&?<:.RV9ICS?LIQ70 
@Q]R"6I>8TJI/&#M>*HIK9"]%Q-$5E26F"V)7<-I.(14 
@<@*+CL\/7DC]+^#(;<@A,8NW&]-&W.U!WG>IH!%5H,T 
@DQ%'>K3:E43 $>? DPJ-^?3\1L,TB3$X\:N2KNTVH*P 
@YP&B058EW4 ^]!5IOKL>CI$F)"6+Y5C#1LI4193>.(L 
@W(UPUT7[[1%1/1LMH+_:>CG"B^SI_FP.F<FR <PN>$T 
@R(\!^:V>Q]_.[*5T-$'E[P/B _Y'DD+:\^L2]<8,*68 
@NFH+9%]OE'*(V%K.Q&[BG[#)-DIS%9!6P.$(J7YT03\ 
@?WCP\.-]O$XPNY+"$KH^_F+5TA50::X;B;=T]G1S,18 
@+BY",[E_*T\"=V@^^@_S#>9O/12#4*26B0>,<'SJ3X4 
@9-S];TSR5KD 7#)KCPH'O;=?YRUN);%O%5U#KG:_.E( 
@SK9],"UEC:@F@&31I\(;AWF]VH-3:.NI4NHY(UY>0[, 
@S^7I)/D4B_3ZVLZRVXVP'<;\ O&5.4^48\#I8SM*;_L 
@=8I-1L44G5YM!05"&U3<638.NF- S$' B>8V+^!T N8 
@N#R.5L%MNRPM>>*!(76UBC1ICK2)JR7E!!)-KQM)DV< 
@'Y.IW*2YOU!M]BUX:\"QINK\H+VR4LM!730QB$>TX!L 
@ O=%&\?FCA:QO-7!=2,8</ML?VM\F,Q):MQ<]OH=N2H 
@'>UNR6F-0K"/;][[(Y98PE'!8UN6N,763*',*]Q,%IX 
@7R&81(4W8=ZA(J<^X(9.8(97DI-6BD<^;4M T-_XC6T 
@VJ\!L>&TED'KEW_"NH:30#<*QQ.6HD-R#(-,4=82J1X 
@]U!6F^3'> S)%P@CZXIP->.:6RTQ5^A5F@?5HB7,;Y< 
@94] 0CFX#K)81#,1*:I/?8V./C@4+<,T_%L[X.2V$^@ 
@4!+F77&6S[0R_=ID =A;3N0$S@)@A>?7Z7;%]LA"V*H 
@9-_,I$<KVHVCK/=WX:?@J4OCK'RQ\$W )[:$XIF!S"8 
@.?DGP^$S=,X$<EWR23>'7[N%@)>HWK,B&:1#<E%8YDL 
@TYES5"0%@6T//"VK)_Q.D@R=-KDMEBC-@4CBF*P8E>, 
@7YL>4M<[+8BI\>GCOFG36F"9=VCRA1&PA-]-&[/R(;, 
@E,U, =4H^]"[4*XCE1^#N$&$C >E5+P?LK![4'956S, 
@$^%XAY.I, '2VK[S(MQ%/](M\0F5613;J(HL,B>4D_8 
@X1XX,<8O'$@7I>'6,XV;]HTT?D1MUK< K'"X$Z/_?^$ 
@%%J"PF\GAA2,V**5HA;?]=N94=("UC;$&E7_3-"7^XX 
@"KP\2"FWD^ N'LV1#/KCUP N?,%>_0[DE.6L7TV_T$4 
@%J8G)<;\16)2=:3-GIZ+8%:DF?USET2"7#VF!0VUH?D 
@<)PT1:.SU8M&(KLWNW+JK<W;<3I;:Y3:QE:MI8-J2V  
@/S"*C&J* X&0Y1JG51%>M]B:)<-61;Y0 X_VE]RK3=L 
@J41V^YH#VH:9H.LWX3R6G*C@P0C5!2I-4($@YFB%3IP 
@,]T]3I%F=@B8DKT8(7&8Z&T@M2Q6"_P]-JO79OKFAFP 
@OQ K2.L)P3B_0<%/F3)-%[IEB2W\QP^P;<;LO':H4Q$ 
@W1H)ZJ6)&ZHW9VB&1V6"A;*Y'.R;8H4^TU'C^:72![8 
@0?(#6!;G%.C<$MH^H5EES_O[=0$YIT_V:<C14N<CP'0 
@A^Y$^:%#(H[RZD?JY1[+W$64.G0*7)_OO@UDV\1^]4( 
@PD8PWFPP^:5[8O3Q,7=L4'5^0R]9QVHG_AL0FJT]26L 
@DOXHP(Q(PF@.'ZA^HS!W[O]BB3C.#J[\J3O(F8W>DRX 
@AHS\34QXE]FQ0&GS(8O(S P9/CS^"2-'>%9F[\6B3T< 
@7N(P./]V-O>6SVY$A71CJO3@ I%5VNSY*HSMB&\6$HL 
@YOSO6,V=^5Q!7KB:#".<L=EV+KUZ)\8M%VI&LTE?GTX 
@I%)FV:6V8_.?= B)8@:IY)9"NG('WS[7(3L8EA<0KYH 
@-H4FVR]]$NC5 SG%FPV?&J)3.-?8K9ZH@=J<;A0I^04 
@W#9LU29U6 BBYG8I0*,[J@?0(3%=]XI<$'!18N%=).D 
@\=-PEK)"H%')@!EY#XB ?S@];U8#2>K/?T]G^EJ(U3$ 
@"B71_^P=-3V='3XJ>AU2:)M9."N2\Q0U>V9&A#LO-74 
@[+27],ZB_,M2\Q]85(**75"3L$UV+Q?G;I=?R*W84%P 
@MHQ53@3 8N3<=3T<"YKWN/5JNT,N@XF!RJ#XB)* PAX 
@IJ< 11A4PDT6C]2;KS'+%!F&L:6#@?G@_FX]V7B9>TT 
@3F 182S:D^'(#+S\L:V0HD>V4-RWZ%5[*"E=CXID+^L 
@<,\\VN$E=0U6T\.*\B.^\Y,5F(D+>QLR";XS"!INE+< 
@-9OQL/.<,!_HP9UO061E%^_&Z+'HQ7UG_YOR6[34=M( 
@9K7)HZ;I<2]=Q%$1#?'@]:-FL?P_9L1, *+ S.QO-;T 
@,72544^SL@]3(8A]017<PD=\]5XM/D4/K'!R)1G";0H 
@&M6=.VWH"NI?XCM5HZL(+KW7OQ)TJ0=>4U9KZ@Q3IV@ 
@/GKQ8GA<,(^N%Z(N#5Y>:ZG0WE,IN(@;PT*I=K_.';  
@ASX W]AO6"'0-H[::5*?E\L J_BJ[OH^>Q>:XY.V;PP 
@[6 $1S;Z._+5;.UHM2ZFB0846$H-))%^/T=T'!OV8Z4 
@E58H @SNI5^>&<@SG!916K(DJ*&#H@+PO,!W*\GS1^  
@G7MF4&DO_7779LQLXJNH]39E2ET[16_]>W>*9C&&R"< 
@=":$8_N)J9&#?%5)T;D=(X?8F.G("K,8]$C-7MCY,Q0 
@1$HPXY^F4/FGI!#3(:XDJ<-/ 0MC_UFXB"BTPX7$6Z( 
@Q(-:J:R/,VDU$7HUNB)<5.WUHBD GCPSP0>9!3*ADAX 
@U6Y],K7BG3&T,6@#8T4R*C5]5?3>/N4-W1$I3@JEXS4 
@!>S_8/'FP+7!&A;660R]A4[NC>QIOLY70$&!'+,!-V\ 
@#0E;J73RRTTI;IJ,(I(PWC6U2YL6JKF(S Z\<R$*LP0 
@B*ZSR[_BI<=N6[EK6V1BEQ%!O;(:L6Z %)VN:6S-7;T 
@&&P%B/9@_/7U:0.D<>UK GS87GM'HBM)4SL(%!"E8)D 
@CBN6XM8X;BF5M@5L#WZ]]= WE+[X%O>PH-PZF"WG9'< 
@K7=Q=92Z2F[#RYICWRA6U,.:?![ +J PZ D;\BH)#+L 
@98%/B1RS,1#ZEZF?BRL8[+ Y:_P.,KO,W[F_7GW-9B0 
@R_8Z.Q?1F-8ZN%AI@2])IVYS4S\BSK</P=ACH22U254 
@\9).LI?JO"&#Y5$LLY0&1C.BB<GVN!6*%Z-)AR%6]@T 
@(0)!(DD#0,>Q498=7=ZI+<:O#<\P3ZTBNNB-O+C3YU  
@!!8QPUJ23'0/8LDH<*9M>'P5O\X.&](2!"JE0#7AY*< 
@Z\M/?+M.8]H FY Y"8]FNQXZYK76R&/AK/YS3R I)/< 
@$Q+K8$=1]$#,<,X<(,2&'XC7G9;2H9.L31;0SX6.URT 
@<S&PK,O1D,_MCA+\DD6;QR7+$7 J+AF@/[3F7B^>E:T 
@ZUUTW81\W.G5A7HK70W20M6UW><JI_4B0Z-:<-<YYE4 
@7OY@I)GK3LF\:EP;X$;O)DERK?Y2BDO!74_<S.2G5=H 
@Q*#$KHG9L=]MFJ*(JP-!NCL2 :<W<48Z9%R:#^YTP_4 
@]\SWN$R5@*EWV%*>JTR_/@KB@E0W'Y'V99&:1:#I>^  
@A1\AB)-D@+$8"I96A>,(062+=8PQ3QZ;J$.?LJ5QLB( 
@9H@18**<OP&1J,4*,E9-I0#9\O*LYITVAZVXONZI]+$ 
@_&HMU;FN<37"G57X8DJ(]PWQ*O]EI?G0"X5%SV::OJ< 
@7N^HW#J3QZ(GC;&%RV(#TUT3:8X=0?/$AUSCJ;4BA?H 
@+6N5T)(!F,""E\Z2.T"E 9%=^^4'E6U8TNKK?;2]>)\ 
@$0Q,P\4N-\,\E5Y0)?%_O=;#;<M>:X-4 N<$.XC.']< 
@%A40>5-MD\*M[L\.^$X8SRCAA*3;MI&N45;NU6 6J-\ 
@B>"!HV:^)F&><#H7EJSO"[!2C'%AZF?G7/;B.,K)'D8 
@62,NUG;I2;:F\'O<3WKPN'U$$3D!=-)211MG$(BS9/, 
@0>27J:L&,=2YT665]JTUQ*R%I;8F_.[+PG.]$Y9USW\ 
@V-P/JF"4)%(%^+&1^C+,G18V<LGP=J5,7/?"WF@&[@L 
@IYU;:]"P #ENWN?]&#7](=F%1J@#&$PQ.)M2*]M3NC, 
@^(R<X<>5!CD:A>,_E]>*8S9!K1XB.T7I/O;$>(Q^BI( 
@KTLPG'^@%@8VQS'CST<(?)EMXWOY;12L$;%1$S!J- @ 
@ :)C!QJ6USRE8Y8/+P"<L-'*PQXTY$GKJV9;\W>"5-D 
@B-N!Z_(W+<YFJ>X\N U5 A'4UM/%NK#0/44BIB649)L 
@:KZ"*\T9WI43(0Q,<T=S4<OAV06-%%S=1:I;G?6+,'T 
@;0B :+*$$!A1UE8J)ZV-%;B]T"Z0119'#_;P4=@3&"@ 
@B4T[2D"P(9 */29A^%.O9T,#"NG0]U7F^" T12V,0*$ 
@U7.2ZX$5EIOL[HMJZIOP=X)Y?3<R7D A>\Q'4S&5/VD 
@ I//9SXW"-6R4IJ1Q2[.OD+=  #,#X>DO]/:APUUMUT 
@\<Q6%W\F9)?L]-(A(,ZOHLDI>;6)>#,G\YI!.?)EF=4 
@92103FA+0Q=N-X,R:!W]=C&"^<FP(",.=Q7)WCIT]>8 
@*O.\?LU= Q(JX.AY_B;FAV<\ <! > R)T)ASAHT YGX 
@X#T=CH7[T.LHQW?6>WJC Y+9#9[C!Q"B*?&42X.6S2T 
@925[RR5!!.VY0;W<[[&?_I_P2OB2F ##DF0SU1H1TK, 
@N*PQY<OYE+\J(2Q .G_DC71X+6'08<6;&(5A2:&Y@:D 
@(0;=$6O**WJ*-N0 YGPW[:1A)/XXJY_$F.^R#5(W5C8 
@5K<?\-L&4SJHF3]49BF>YQ[YCTK_03^Y/Y\SAQZ0CG@ 
@&Q)[[N(>%0\Q-PT\S=]3CZJ8F:EZ)-KMQB.TW7-*3MD 
@1A*"H?(47,,6\JJAX$AZQ<J%JP.;J/P$'.>X?-/B$?  
@L6C+5OA3<JW,9HIU5TTB>P6)J7WL$O 5L6S7=!1I_NL 
@Z@AYCD]J,7 ?,_"8@0NJA']T9)/>FH\>NC=7@.*>/ 4 
@@.; IK-TTYJDQP4*DLBGGF3)G>%0HS D^^VS0Y-J2BH 
@UXC-/>A9*G+\D67#_6D$W1?P#4@K'=HX5H-OY258.3< 
@KQ<5?$;Y81 O<:2*.YQ+**S2S<=P7:_RGALH\&#^9J\ 
@8X?XRE>L15:R)6_,?+""?AQG%A3BH('@=]OCBN]@.C< 
@0EKMZ/^5S&?X\Y;LU,WRUNLL,K\K#I'4N'RFYA1A"L  
@X+5@%:#P+3>+QAJI758QTI!_Y,*T$C5Z5]$$1/H[ZHP 
@!P*'FNM0;8E3A0@15S*Y+LYC$!#3WDPJS,W)1E")2JP 
@SEV5:!+@NH&B>,JC<Z%127JD]Y<,A;_Q%EMQWO]J,:X 
@8/TK)UHH!R?\_:23_,G!1D"V=K8N;P"08Y2;0?+G&9@ 
@5"*(@!"Z\/.2E5>VK48R?_HXC(!?L%KHO,F5\:[;*ZT 
@%N+C@V;-+2EV0'UN32#/1>82I_<6*"R;24B: +_1.:4 
@YUZ8'C%"W[?YN1Q%#JVTS3LX3DH?2\;9%;:Y:B)%<A8 
@0R2LA4U3[,?!:>;P^,I(*Z#%]_5NJP('3QA&NW5M;L4 
@N]UR,,)-53CJ7,R:9"$J],;E;X?BS"&LG@J<R2OK>C( 
@HOI@?Z\Y'!*CA7M'(Q+_?O++XKHZVM?4.*LYUQ /IQ, 
@-$9%H'#V\G$V*#)9:G2_)<G6*!Z.VCXM>KLC,LBR79( 
@IP*E8.A]J2$@MPA.J9+;^2$QN>\$94:!&PZH!ZLY9RH 
@^8,M6DOS*BHAE11S]T>-I@6C&_<Y0!17RHQ)=DASM4< 
@G+Q+\9H<,6/=NZC,5$Z:=XD3'!&#<!W(/"QV:U\#S0$ 
@/6DQ$>&PUO'L$ ;U<0'$MX]XX0?IA(2WTGGF]KHQL T 
@JVH8/1Q-:ZT;-O+_1>D)H#0B4)QLVIH8396 B $T16$ 
@Q(TU8)C]R=XDQU$86[6[KEM8H (@@MDNEG9GS&4<+L8 
@W(,4.J)-"KO$SSO86(R0NDT ;=Y^S= "6ZI.(M%4IY, 
@DX82TZSC03,070E')+32MOS [R&MO4WR&XD(#!VF'?X 
@'IL1^U58SM*?PG+-42%"U#Z4(*E4K"I"$FC#NFWK;\< 
@6-+.ZEUE3Z<7*V!%-Y#*:>K@I6R<!XH?Y>!;VK3[\V8 
@"DMF-N7PEM(@[.+F.*9+FH%A=RYG8@X)BW^/;C,4OO@ 
@NU.>47<H9*7\Z! =#QSM'VNNB0] @0K(,%.Y<Y=K-0H 
@B3@/&G7@6"N6_W^& ^/O J&3&4]Z'''Q\V$J?Y,Y7MH 
@\?*1>&NW+K&).$'*# M(R/FSK'8!ZA\FDS&BE@'1"48 
@O?C*([JZ/7YHGIJI%UUY_^F\@WU7UXCL\I70#39POK4 
@AQH!0Q0;5 R#@>J'\S%/6-^CT!K]6WQ+PW2'0J6)H/0 
@U>K.P7NB,UC6:\3WH7$^2FLL;.=D3&L&K*FQ9(E;2KX 
@\E9MCBPB,YL+B=MZ$W"Y:O]>:1%;8RMIM2JD5IG<O5, 
@S,SSQ=358H8WP:'6)(/>QEL  KN$PDJB\8N\ZP3.#]D 
@M+,)EAO/&$D/.,><T*!6D)U T+FVLA-?2_M#,:7;+^H 
@2F4KS7L-)B0GM7\156L>^7)C.IB\*^C(ZU^J_'_S_4L 
@3FZ>/QQ L4B R,_]PI(F1HX_7'"9RA%4WY;+8]4UL6T 
@?=GN$ZOASGG_J)!.UPQR49OP\5T!8HK$F1P!G#9I/>< 
@6PU]V?7YVR +4'G*( D&\7PG*\'[V_MT6<"2](@!.>L 
@3U=FX>_&-GRI]K"Y?\=H95?;2@PULT$[)K$A&C5R-5P 
@R@C?C/=OU^O/0LOYLH =!(5D,.WJ^$99X^!F[M/87S, 
@%??&@B$U9KIVPYK5:HH<T@SS43NW^W#4$+_5-S&;%$X 
@/>'9W;7P?W\?>J&O+[&B>I'00I]5U YH%C/S-(H+U0T 
@KM97$DGH\^3<CMS6+MY "\UX^GFL<A6V15,3<K/@KWD 
@_3T?MA(2\6PL/X;,IQ3T^[@P;W&+\;I_R0#:B3N?U>L 
@2[D%.9;GW-7:2>J)_0>XA)9JK;/&J+E&[=9.E=^[DTP 
@@[= L05Z_1ZYI'G=I9(J:9G$VRUIQ4G;.K=[PY=A@\X 
@:(,K(,6+Q+301-J9!, NMCKQXQ8JGZ0#_F6QW'8XPL\ 
@84%Y*U-43@Z622\I\)>:9<&.BEI5BM,F;FHG6D-5-G@ 
@TE=O::"2YT(O5  K3)2=EE%A,[=\_:"V*Y:A1KE'C#D 
@Q9(6.-8>V]7:8Y(Y+_IM/3&.SX,]_S;<-?Z'<,2)PJ4 
@VV?L\'7O 6O<TO#:>#'92[0"3=)@76NP/%,E(_H_$)8 
@U%^@#U$P.DI!M;]JS6#]GFKB'K_DE0.GJU4F'&UVWQX 
@],Q'.I R9LK5+)0@IM(*G(;]$,D0G!-^+?- KR5BD$( 
@X&V</5VS"@TKDL")=<Z+U%K0U,.MO:YY0H #IN(_LUX 
@C4Q'9AAZEL9LJ7CQ,+7I7^?$D# 1;I*FP>]QMI86^#4 
@H*,2ML,(%T3<<EAVX@3MHXK\=K(7+$J=A\!HP&D&H(, 
@U@LV@NJ#[?YJ?PIAD>JW#WC-/8.9[XQ%5@%UHODN\Q  
@;T,U4-79#8L(94/TD(?'4V.TV'10/*4'>,+Q'X%D:6< 
@NB+86Z%-GDP;]> DLY!E%RLV+[R(])!)VK_N7HHVF7( 
@H=CK4:[Q7 05P1/CR3X0%=\YXD#S#,5<&Y2&45* (J4 
@#Z7>&Z84& ,JL=410\]W@NS#EI)I(49EW7O4F:%A (\ 
@;_$B7>0(<,(Y;':>C3O,C>SY;PF]US0>Y,1MN>N<0'\ 
@@,"/+T"ZR)ZQ:THC((:L+E7(!*,9'M(?*MG<=S8.;V< 
@%<W_6G*[/)-:A5US9TS(R:A!MV*!G+YPP+^-LFQ+*Y8 
@$5U.WB_?)-%<LPF9^=?6H]Q *T-ET3)Z 0%YMC3O_4  
@MGE;\2:$?.@=V4!H%SF&<HD#V0;#(63F?FG6V3DY6*D 
@<\5DC_(JG92NH3P7S.='1<Q7<O':AN!NQ%)W1O@@MRT 
@XFH9/;])4ZVVBR[U-=^TGZSS #W 2*E_]_HZ,()ZGU$ 
@TC"D% :U1J,4E*8T[(<Q5+$JJ:3Z*<NJ9N&3FBPLS4$ 
@%T^-HEB%8]HA=,><\PKCYI2S%IIJW"!GF(/IPAJG;XD 
@T#'PG1OS,:7QP)>Y!52RCFAU PBE \0[+;@XX<FXZ;< 
@_'FH+K9:&V!@M^I8R4Z<;_)=3SKST'ZV!8RS8'HIB08 
@MT^C1^4U-I+E$>SD5O%KX;^I]?D9Z1,0MFRN()NS63$ 
@6%NJ,G.>(5!GAJ9#^ZUFN@< ,VE)0OVA@;:2[VM<7I< 
@W36.>V%'S@E\ KP9JPE\R_]YHYV>\>TG,)=6[U*>BO8 
@S&,MB5E2!*(MY IQ)0DG)=G#/Y3SS=.A\:8X.+0Y2B( 
@=%-AV !2FL4->>HC$NSQ"9MS DC^CTHMF<%\CZ6K[Y4 
@AL-HE"TZS1,>TRF=.T;[2F"I QZHJ"ZP-/FU!:B#!4< 
@)*INN[N<,:K_Q9&Z@HAN%,_C,-X3B#NWA(1I"]0)ETT 
@!]H=&-?4OUJ 4$4OM]0MOSI)"CFW$-Q.,H[V5!UGU%D 
@7=3>,V!T<66UE$SO8PS J_LJ '^U6SR91<"LS^#0^P< 
@Z:P^CDJ*9I[)D_=U4ZVR,]0^.M[_[</,]A[DJE8U9>< 
@YA&9[Z<4;:R/\&>@/E&^YS\UE3_7J,?HF^KU=>4?A(P 
@L8<N>&G$LR65@7"'JENC.00II*;@=<Q>'H!>#_TU*WD 
@2DWJ&KQ<Y=8[-99(^EEI1/"M(IK=P ,']'0RX\-(YO< 
@A?XZA21[E_OJT+0-S<D \5GU<V-D/CXZ\&/-%(6^W2\ 
0S 6X"W3F/B5*MQD059=.#0  
`pragma protect end_protected
