// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
J7snypruvQiSSvgtvC4nLt+Jzqex2dkCwjWz2s1at7OfsR40D1NVAbhA3+zdd8+ekqjU7eeDfpza
IRw4u68U+6fg4htjLbVV/QiMu7/5rYAjCjbGs/ReTTZx/XnJV4rgDoCFOnAJsS3xf55Fzq4KObsv
brQMj6xT4GIZbd3mO6/PDnHStogADbbS5YB7Gwqv+mbgpGTGh6SkPdjdUd8vfqKev45Xc1/7SY4q
hJmpWvfbtDC+fuGeG8hatsH1e21MYu6iB5DqmUOtRF/25RXBr6WG+z3DDuVTkvT/xe8nqbUoekpq
9/Zi+LmvMQIAIS25ZsSe4I46TNVb88rsPS6jlA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
yjfvRoaBEpCF7hXNu/H3BH4FIGHd0N7+LtYCGXe8l1FZ/Sy8p2i2UeTHKr2iI9c+inr6t3Vihgh7
4BC/GHh3xXPcL5Dk4reH2XxviTooN7cbrWJJ7E8TeG/8wKK+WMKZEDx5i7y7woKzqASGJAQeADCb
4/ACFhkw1GbnHuCoWzK+Jcy6C88FyukOWnzuHHUnnY/KDvVn16M+ibkJTYstFHmyR5v3MUj1w0PV
e5fPmkxwAbwQ3njL3hWWd3gWhnoHHcLbvFQXvv7zW3teaXPA9U2SIQHisSuUi9aeLnqgK5hZqfyJ
hoj9Xip+iTqhi0HZBAYCBaEr7Hfe36cZQJATfzQGgyUW1scOuYbTsaDF+Lb8+iaZDGh9O/raw764
2/awbNIxdwJrvZvUjgO3Kh4RDm0w9xw3BXR2PNHIYDppo422zY50IZJ3WwUEflydo1dgKDg34P69
JRwGsP3ERN/cQq5kpdA6BFUcbLvpEyNN3O81sQTiVdUgAMUNMdkMbh7uiNSmu6cy4ACOT293Y3vX
zDESOwGAecSpv88uA9AKxMiL+BXh4/ZITY0cmjh7oRq401r331X6+lFfkyZTemV1gyFo1kjVo6vf
clVzbKVvmKAmDzdnHPpEmt3qFAqHgwGUD4eF6H3sKppQG+TbJubDvCOlPttZPj1LgPus6IqmhcvK
g/+GwpJWtRSBgvp8ns9MtnGBtLX/tNTxdO363MKS8daN4EeTdcn2kTKfZwBYTFrxag9XiN/6C5G3
z6w7fAS4ttaFUFReGOdy7jGBhWAvrgLUWjHUtlCk1JU3hawJALAMsntWGJLEhsqU2Izt8n+kxPfJ
p7GzX6WwPfZCX/YZPwR2/ARrLRVOX9TOLvqLrNyGHEjMOK4Lsk7L+8NLi/8/PlqnY0LFRVJbsa2V
1nExMv5w3lAAnmPYNq8CMBnpqv+V8f54/wR46vE4qD6+Ek5teryxcljINSv8D80h4JZT6EjL2pSB
Iit73YFTkBcXFyu0HFvEJWMxtBZ8T6/qsNIdKSI686dIkozgutwvpf2rOwP6jhhmcYEVNd7gF/Ra
9zNXLcgpT692Bwrf3AUV3fXkxvkX09RimFKfd0P2igRDKiBnX3fvxdCwIBvAlfqzA/m5G5sJQF5U
L3hOGZ0dJSQnEoKgAcQrcBKQHUvwtLFS0WjSn5hKvhtZYBvpsSFkE5CznImAnzLbH0DwzKxNv/2M
I+BvMT3XVnctGYD2ZMvOjcPosodcM337Qg6i1ebim2qzJAdSV7TP+Ab4tDLo480mA2QLIdu6P/8V
v4hvC/ygEcFz8NvgwVzeHD6mwekNQBsl7/DmhCP1XdYlyHXvyr6GEXTjaUoHH/XK7GGoKsJeZM7e
YGaaT5omZKUzze2/8e/vGZ+/Tf53rNHmubNY8vU7j513ApZ4qfCVutnFXHPp7NoFbgt3aIQqQmh8
svTOLDVcdPPdTR+LWnz6NB7Yy9tR/TQzzpUEL9vujMHJGLH95ymMfnhEKXBtR+SBFuahbIsOu856
mburW1I8o32QIZmrALaztIOjGN5fqc0wHrDRo1jHeS6jNBUppezOZMDudZSkCvfSxV615bhdPSRS
64VvxK/NzoUzl3BJcu2FXjGl8gESIG0ywxA/+DikRoVbwwHzXYGwWKI2Ylee6k9oKi+BhljrjDKC
JfoT72NKFZl6SFJrnc0MWA6csoWJLymcEsaW6m3+pWyT9TkpV4rwvDuYCaURYmMthKaZyRjhG403
++8L+TkvKvaT7WmOKFmYiRae0Uhm5UjErzKAhC01YX4aeG5+ThV7UiyUq2geFw9Gj3RHOQ7N1j3i
EaYb8cnv4f/hSDxW3ePZMjF2kyo16sUebBvj4mADnmDhcu1ZRqPnIVLCz2CsacMtJ9EWqopAt8G7
el/UQpQNiNjE5i6nXP3CyAJfOD9PJolp4Pl6M2A/QUqpScw33VPN1EgH0ugaYZQv1+jeVeoTWTK4
k/QFbjfko/GO3/khsw4/05lXqHu5nUBvshBXNVomaf+y/FRaryBFWS3NbXG8BucFiwYny7pPaIF7
Ey2Y3mkRjMqWltTrRY8/B1KOXT2584PdRq7tE4aDWtz4zkQYttddG7pI28jRjJhiekUZKFlC2wLe
5VhNhlM1oePWgWiIaZhqL4NWrHJV7ccQSuCy/2i2s7AkWQ/Koq5nOYbRcy3yYQiomtJL/nX6QIVD
+xNjViTi1vwEA+LQw1uZa3hg08+XxFNos4k7+G8jBmn3LXe2ODsszO4JEiEnXWjcgG8krx8pdpjA
OLwV5pCNXOBNCWQVgheK/BGyn0QDdti1C26NSjfg7qjkvrxRf37uTj24+71qvKIKawvZoh9g64bp
ebxYTd7J+wzInX/BZs4EkhzV2nFjCFmfAa8kjx8kztW/9SxA34vOTmemYT4choq6Lv3mUy1GeCcH
jP4Ts8jhUPfgCGdSuiqxbGxyonhTQ9Du2bJQ+LRDRgLkkEZen1C38VNY/A6/IyXrpMnS9sMnanHR
XCe1LtwKqeAM4cqKDbBZvkqZk/vqtEtlR7B7KxtsLfqe2z6BxgpP/4pOq2tZbk9r0QgSz1zqZz/1
9DD9UubpoaTPVF2XXzAmSK2TE4AehKuvr1rxRawFKuMbDWuYbzNvlYDdpAUHY2WRp44rvofakzXQ
g4cVpfniS0krrgLE4PmPdlgsnio43f607UyFtKdfXovJEhLdHyKIwixAfPS1tuDRZEmBOw/I961i
yMXOr19v3RjKMbIFQkiBthKwQhaGYlw+IlKLvOLTmv1kGU7HjjYGP9R+mCvWiYS8ik1mR5lJc+sA
smW62Zn6MwyFsVnw9yCpH2EWieZ4Q+fhJnEGJgJKKd5IkBHa//0yKxjeSpxQgoVFY9i6UVB3mJ+n
kkFgodaMRz5+pMUeirM7CRFyZf0nNvtzf40QOcQtoBP92FtcU5QGyE1/htYMVCm60exLGU7XPbdQ
pRAn3jAu6r2iB/4XDOst1WwLwXfkX7do+UBhYI6QwXKAWIKjEG3ASB6WspmRb1UHv47cPaGhazzM
+LYJhqQRmeADZwoHkJVBRXag0i+UGkQFuOQ1OjwiPnrvIenqnafOT2ao4PoDFo+pvH8l0XPYaqJq
Co+NxtU5NpdoFqxwgC3JsXuCzG9I0NzO3wEMicQHNuxg1WofNr/+W3mFTUARYZpODBzkBd11AaFx
/TnaBp91k7iz1owgtn6ui0810HL1KSJBcCv92DOl6LUqoaTQnjcHkVyXJNPHKkpablNusE4osiV5
0hyTd0viTkYaufSfI6IiLYMHw/KZ6NPuQK1w6C37PdHDVVCYIBeLrrYZJoonYk/1qsALXKjoorlQ
tKsCUPLO+ZO8MDcNin1ATrK3zDGqIXNByzk/T++aRIs48vfUGykka6IdyxemFDKAhgFMZA4qawhk
JESgY30l5Ql0BAdb211HajackpLEyGmanbyPLy+p7F0TsasD/l8nrbLXe1NBG0Cuiw3bCbo8WAZs
JiGcF8b4EKyolTssnaL+yTAu4f7DiGPpU8Axhw6TYCKnx0RyGuuNjWy1ZPiktNygH0M+H/puW2Fh
ZCufFy8tc4R+lgzlBQjtHdi7e1IMykv6YAuo3iGTOuRDtotnoVzec0hfJ8Q0XZiJonsjc1KBPWmF
syMQonECOmu5q90Nrm0I9BQ8u8bq1afAuz5opDLwVgHc3suJYHSTPYYqwqDjbrQQMz8rgjSC+125
/GI5g3+Vtmsrd5NHRQMA6ehKwil+SVZgZKwwmD98KsKNb3PRWdx3dasFCUHl/xXI50oADMk1C2N0
c79XEHBk7k6InxmOFHXuzl+6PmCWa3Q2iIoVOH2gMH53CbFBaO2DgQwcAShJz+NBf4TndHShXd6j
ngZQH+p7X6JomzsK1IfTDzovtaJKr4f1oCjs8zkOdG2ml1x6MzGtdY+ee5crsoa8g1Vi72cvL3Zp
Hkp98RsJX21IFoQkflcS7CDI+DwRooKW3mo+OivxDQcUPW/8ZBt33ZjA6OKARS2nqF5HKeqt1gUm
Ueknuo6CO//0W/4HGGN929SwiksCfK1xDICb5HZ5hmz2mLuJZ/TrRryQJtcsiDc6X1XnGYh0XU0G
cImXE1aBs6qkTRSNTIWOiHXIwKOopEnYVQRo+jG0vcloXadEPcdOLk8DyiU0jCLMY+LxAcV6oDaS
jSlWni4WRUFv8pESSvh0VLTE+rtTetVXA5ZpGkiT9G7Xeb/so0iSM2KEmoS9Po4C8oT5oEWivGbO
GT3VmBg/g/7Vsw7qQtRYLBl2gJrMjUs0Zj4Qbl5rK1kqm81Ekml1bf76wXHpgrsNZl+wP8bP2TFk
TdgNqMyPjlpxJ3vm1g9/+MD9JLZaAkHmSierLF1dAVtFzPJZMrnxquju0eG3g0ravSfHBI3c9L/V
M9XQv9ibVHc6LAcPqft+ftNqZHF3dEOWrkxDIu4EVy6iw8X8/zh7xMBYK1p+pxgREKSWgXnFPm9+
w1CdLucR3Hnv1GR7ZvKUrEiG/Skciy8rGrgMm6/uyUb7xyizPmaQ6bNpmwOYcn4Qp7/lK+Oc6tK3
a4sd8HdofrRB0rF5M+biKMHc22jupEjfocT+jNXrBqQdGycxtkGoi5tG85hUAOzAURVBp3gcbGQw
kCAjgCYDHNiTXEilTzyPAsV/C0Znhw74VqUFQzTBLJ4fM58bq1Z0XrxicqW8VuOWtruq+v0dSfui
YAuqIXCJi28jeDxEdKpMIfb8jvAV9X2PS4Bov5j5/ot+ixt/10q9Mz+YZQp66AdsKT1UIuBoXJO6
AJoskEqUZer0/VHiTR1c6m1lQqAskRM2qW24AzfZ4qwQtjRWFCs2cpw9M7kFHXCoQyDDqKkheVd9
0I4hCPSTbPgj+LV4d3BfzBhAyJVsaalwVmGus2UMLEOgQNoVHt6qmdgGtCcMMtdFoEgE/+STkxw+
YvtY9ZOdm8Pwj++4UUt/zQ9rMwewyBhB3p5Tng51/eq0kNefeUzQQ4+Z7LHy/4gjuMeo7740mYH9
3Mw0bhOUlWnjP0gOozqPJnyjD75Z9cdUVTSKwMy7jBxcU9j2b7PeOwNbPUZta2TwBd8ScUOplBwz
MV93PORQdzM0VR1FauuaImOk69akLDNnxTsfkmwuDI8Y7SYSCBf1Ay6wChigm4SO8gymrCyZnYtA
pddbygXrWBcldGpUp75eE841zdZGMc0JyA6E4nnSYhLIt943xZqa6NQX9QZuJfkQRvFvgMSQEqdh
YV7tLwqfhGk3LRSnz1ZSWBug1Q06HDVd4VCx2cp1KugK84UVaOn5AOulHA0lxiQNoDDJhUb5FHh2
/jO1HpYk+5J/KyTW5BBaCbeyxXo2HMjJefwihXOPSOC+KaE5JqkGr7YZfoWUjQJG17Y3u4VeJ2fe
6pLmknL/m02xe3QM+3GowuAaUQd2t2NO4I0g/F8vH9Pz56YoyPvCFB8ZcJC1tfG1ojv7H/wNsA4a
NlhbFfabtWaOZOoE97uWi6McKVSHxDdYFJY7RgsFkBq7QeZDXIMlaAUm8gWkFOL4RneNHOio/NM8
VbKFV8WIOLCi4Ycor57m7TVykuDn1AX2T6AhGE29WnrqaQptnNPYMrprfxO4VjlFcDaJTMasT3um
lZgUFsmXQa0hhi18yObH1F7UZAR6QEAlgFyCCV104sIe6JiZOw/BChxWM02z6YzD+PxFFHHG6/3l
6rf0VF1FnQbYeD7Iy0ATvc7CoB/bJpoRLsisnVM7nuW0PdyHhyu0O6yW34viekG+vQuDmyadXJdG
2+gb1KOCs1G97spGwH0APdeyLoPxEsXoi30D1NiXyHetOXcaN55G8Rek9OKzLmfYRWoRufhKx+JI
3M7IZPQr06ZXya34ngD3tWnZBMbp6jXp3VL6brT0CJQkBvoBlYhNAUf75mdzHN57A0zpCRBrrkjf
nEa4wNIITMT77Ydwll5WZ2jg2ED8wcxrw2W8E7Ih7R5a6oidIZqHQEe8II4782S0Ea3OE+3gOw2T
nz6hEFU1g4tyEVr1+AqBxDxHD7+WnBjf1bj/t7tYtvq/dK7mgNnZWa/9VSTAuA0fAYAIT2ON3vMl
yHaYK0t9duuv4nfax8cEXRjSiz02qB2pB8cQ7e710hsd5NODYUklc6WHyZ5BurCPOd525hyKYb9p
mcEMySXhmxeLtg+8nIfIC9lCZrvJaKnUTGqUXYqhmqF5b6Cok5DGmexCcfHSkZ8u2p9iGYoOQj1E
SxJRnIjlW2cADo6QapGZlCPs0IutQPspsx6XR0OFxsejl8RsLLKqLdcP9QJNmad4WT4mMnQMKnRb
21xiO4lQwVluRYv+XylR5PX2oCtaK0VgU16PHhGLhaHJtc7JMeT6KR9EYQ66RiMh5F0wtbfH4fPy
lL4eTNxHDGjmGshXLKiuVOEho16atrStRc9D5m3pvcC2wLczfxAuugG7e776L2aNf7c425qBxo5E
FPMtuiuhT6jG78IZ250g+g9EWsrFkBjQ+PX9ND0tT1rjKTZiYsvAePJNoZiG4oW2KG03shyTS+Oz
9univ+M+UNpKR65fhAiEQf7igP3HhsQRPI4FKyGFTO92ylMkaQzq9Cy45flGvzvdViAAD94I4zai
X7L62fLz4lAeVF4tYGSdNDhSpdNvcQQZL4vaTogLM43XljQDxSY6KtJHYeL2UxpH9Sj49bMcKTDf
cRfxqUupYNBc9A7D94pa+HJaLxVJHW/LAcmY9V3giQg1ZIH1wHGkKWe4vSDzUPlStXR5fwMliTVB
wGrNFyMNwZSfSfymX1fVyWa9LhMTXhKsgVPBRdqtD98BKpuvWiYMYhpqTmqOppHabktQQYlfWhIH
yoNj0KzkspjrFTjZyreeY+a5ZGFiYJaILYi7zAq6+88qt5QzItDPglkbtgc9yf5oZ8D3xEaLkFKP
KhwGZ4y41IoWRme7uiYodwHQpglTDhFBRmKtdps9X58JcxIGZzFih8r+9K14nxx64bPNPq0oX1dT
7ZjvEAufgBJ0Kpcb2ExVHz+hPTBIc8n/jRUu8BlxEoe2XD90ZcPu8xdwkIicdqOwj6bfsomrIjSm
+RQU8m0o/TR2uW9ZQu7LD873GBGNzurF+P23Flz5d+ioVx5dLYJHLUt9ygWy4UH5wMSDyuJam301
+ubW4DtJV6vlo0bGEYkEZ1JeXlTV7rYYcLfl6xt2Df1AAg5F88izR062t7Y5yBQVapD8Xa0rQG4t
LmxY0AP9QRJABtAw62mfzGCK5oKjIgadHQd6JUYucSfhdjuVYXa8q1sNB3uIWQDTTovq6GTQi4h9
VtIE/hEZfZOmFtzVzBRCnbo31x2qk9jWamYyQliPscr9nvfkh7141DhD+vvDO8KfDkPiMWnaYLqs
USudWYE8vQS4WkehJviofvbyNpMfukrSqSHPu+JdcecvbO0uv9sK/jpdJNNdKLwh5kRqX4Iu3p3l
i6nzDkYE82awfINupXcUf6KszZm3I8cijPd5B/zFEkNxGMPg0qVVYSYNamJGy0wyAnT5zbZcmr1m
Bpvi4KqS2AUxTqbXRa8rSQjLCQf5YIIE9h4XoEhP4CNIUJ99RvnEMdnJFKj9IlgVyaul9R/wwyhb
Hc4Q5BplelpfiyNUITvNtXuAZfKX4RTfBUf/DcLi/kA+KOxxECkVOA9+Enyeec+l8aIa9gH3DDIh
gj7n8AneFNyIF9Z85ITJBRX4zs74FkygkVNvd8Qvi6EZiQGpz/9OvWGSfFEu5zy+Fv8pBhQE+fPM
4YdWcGopm/6PTYaGz43+HupsZvC9vW3sFa3hmq96azh433A9aUzSgRSrV6LC28cDr5ZqTxGq6GBN
Sw+CmUGPh7OafLGXWJDB8VBbgu17mdFFbI9t3ElennBuEqScEa6HKeWgDpuxLp9yjBfbTTaZ2HaD
ACbFQPhWaNYKy1XXOpwXLx8TIwCUzRchIGfcKL7BSp2+TdVj/fAqEfo4pIxfcTqbVeNp9s2mJBx7
ulBm4cJ5bF3ovASZWpAbkEgYLpO6s+fDAUWWdgzCszBlBG/2sNyxcxEYAWnbzK4/pcETje0hhUZa
qpAw14lRd7uLm5ECdM8lr3Ctb3FyCmupbO1tX3xpYZvyvDTr970UBFkYXnrkaPBz+q2bsnWRRo36
rPuLf+6tDAO1iEP8WwukJzH34QATkYaXMtQtEKY6mKMIICtONvI/5/z4nMRI0IxaRbY0+86Wo58P
stGlakLixRuLloA35X81BJ1u5t91C2dmw+M1PkqWUNrIERZ4UuEBn53OcdJRs1T0Qa4beYTGL8gf
Lji1izTOdUNHaTzDxwTSz4lt1S7FKpMd+ShxoU+6HDaZFeUAFRRu+7e+SAzJ/G2rsx9iCWqx7UdG
wx8NlEJU5Vd/zBZoVdYFSnvELUwcNICng3Yg5uRj1kmObOoBUkqhsbQ1N7l6UHlHRdwXwWGY4Mwx
83T/pPLIGwWI25tL40NaQtcgv5EMZD2OoC1UAnu4KDzcA9g3ojxrmFXr35oRsmxXoU3C7EE5sZaI
qejE0hGtdACKU/fwiZTZAO8ubmrWbB4YfGcl16SZMJLVgTMKaK2km0P7q5Xqz3jjdBgicpaBtFvg
ZpUlgrqtiYKtyDUQFvYqsVq0mpMI58Tc0+WXVbDU0HImsjmnSJFFomWL5HUvzEnk0VDN5yxPSUa2
gwVfLlD56vrebemXHUXSmex7qYgvpykxysJYP6cjL/8Xd/aJL9B3GDWbTjBx6DLN8zfPR6E56NyS
ibPUnCu4d7gwzefTt7nlzQGLkBZnBZ53RuqKV4tOh/9n6HeBmoUZInBlySG1siGf54+7AbM0RZeW
bi5Z1PXFplGXA/Wyp7hjVuMhz+0NPsCPOf5M/OYgYGJuFhyKjP8K18GWz0drPiNELzRn2cvWeoOu
76j/oJyoVTn6TJEMIhPa/HSH1gkYU3NH9Qypk3p8mUOpqAWd1KHDfQr7wJYgqNzovhgzEykD4EF1
XH8G3kW0QqWQ0nZ2zG+6vkUNya82mOOqzre3USa3cttHX51tqGSSSYFsfiGrhDKmjebjexTtlF05
K3x6h7n+c2KFIJuNiMwl2cV4Bal7jICLEOYIzYDPQbK6nhYdW/dn6UETUxtx7IDGu1LD5cjPZ58K
poerIVpyFbNrK4Wo67LNHO+2/sJE4MvIWiVrQEY6Vdb2cvuDhWX0oMMGjAVXljausE+h+MEf9wXx
oruJAnaAwd9GpMxTCPqlIZF40aB4s9l8uj3O4Xnrp0E57P6PoqI0+K1vdmiDe40tYwzqLG3HUciX
yKaMA+xePbiTTqDewG5eQoi5byC21nuRNIO4ojr/l/ipurjfMI7ZFwfRtXDnPeUrUoXYr0OCG/Pn
PTVDg1ZLEMladUKd9dYkKfzu3EPVYg2HpGzJ9zBJEUX1tTWjolZ6UI2JhMzmhZPJmNMUGJwevKpc
Sq69QYCjQQua2exEvxfVuJmFfO8tdvRrguAmv6zGma/zvxQkVTpGK+Oaq0G7ZFNIHOzr9kqrEA69
dl2kfeDyaBNxpWBAfPFor7GkFDXgD+OdeNCSGyf/yEKoF3XLuGW+UwWQxGqVcVTkEqnCUhSXH/+n
C1OpTVPgQiNK7pEnbUwrA4wGPYsikYFqMUjAVfmwpqjaVraxkkik5R6tjOMZ1TEL97KEKqfIFnuY
86IQMSLw7fa4qXlaxrWwLeHLSALTG3FtwJ2ckJ/1uYTZZxuY8mnKvyh4xQxuYZ5AKJB3rdCluvke
3jJmhfk0+bUj9SGHTrynYfvD/WLqvJo9CNK5G4npi0qOOPN9smsaBrGK7Nlf1pVwk7zEIvMBJmOl
DKDXPSLQDCyDdXQK5p8y2GT8QLG428UoyA2ImsRpIYmlHO2lyQf49s45i9F7UZhqZy2ZzgdbSPw7
Fh7eF6/zCjZJ5D+9qZT4LwibuknikmG0kUZE4KqbYEZbjHN+6SdX8IoOpZuwW1hdVC6XyjSnzZ6N
t4rwcss9TfabliQKDVGcDPLk4NfnfkWiRy8mNOMslKmgxgd5VU/zT79iOb6vJaCUePI7e9LCRSJE
1SIwPfhI3s8n/qM6awVuMUnCnzq0p+KlOEpw2D49V7A51GFC5E0/ZT2rgQNljX8VtPMzQouKFGl6
E2+jiZmDvyYa7noD88dOpQmda7EOlMTE4QSqcvNNTp2BNtGgojcrCItCwUe/Fngz5a8ZLKCRRn74
4DyRegtHGTI4Z/goTxDsXIItoSuANxIl6t/hXTSwLTKFd5z8k+9K2HRHL4zIB0kOFRxeAA8tCXFc
3eMFWZZaqADDac+/XWNMzpsaKX6ykIufM+2FJKSg0qslMvLgh+V6YYa36M9EI/S0MJtdrpCt/ixd
m1WovZ6WZLY5FEEuxEF+JLLbdvpGb9zoLYIChadN/mG0BNwJG2AzA4UyMFKOcPogMiDAQiYw9Fn0
DtCeVndugA1I4CVCxr64O82Sg/UgpWCWYrBzDu9fok46I15XIrzfyOx8bVnaCQURZek/vrjIPB0I
y078tawO+urH3cPN9OH1ixXs0QBGul2xNo+sWkUnSWD51rmdYA0kNAbSZKwNLEBV8Pn8BZIEkUJR
aYCIx0OKal/ITCzN5U95dQCZqmplZI+Sy/3IyvqKFDhobr52IGo7F5eqbz4m19eR8QCbzn0aAdjC
Qx88jfhcCCGr9Lm4RFB2SDozwSWkpG3t3yg3etYJwr+gpsaqUlOt1fv8m4kFEtrbtYtYe0UlI4Md
Ps5po17dUHc3M+2iPj3RcW70svqZ6JP9kspJnBsivaYPCUqwMO6ZHpqXuKf9RRDTMpKm/YAU1Hcz
Io3pyuVukqQ4CP8pYHWxdJbcPsC7CPhAD28Ya6rc/pzEFZ7oPqj30HMfIvCAEzOhCkEbjBvK9YFW
jznuktVZBPHQ6KrS2/Q19H+p9AQjLjDuzKOZqPYTUn3HgFUUuNRCPV8TERBToCPFPJ6yYJz7OWUc
THsFLkrobwXjofTh9oycS+6EkMo096eh6SdRrNy/e74YtYqhhZAaeFJ7gAmCoR22VV3LKUEMDIUp
UQS1jVvOvs1i8cHGWg162TByFBOQF/7ZWwd0MYyxhXqmq9wjtLm+zhbmlK2oX6uiOFQFCFnN5EXc
vb6j3tPDkSnseTw47L9Jhm64O3iRwcbX+7dM1c4LsBZT7ViBqSm96So9XC+XL8ueduuKzoBqB0VB
F2xUzeJG2KNwjH8DJ0hYTqZZwLpAl8bg55heHAnsK9L9piId6Jn4JSLR4vQk08fFtmyK6xWMIkpT
yPHfltCA4eBMPcGOTNVqG7j28L5R+RQPzF+zA0hJwNgXj6HRscBdXHqMLpF+SHDRd/hBfT/xNi84
+02+aM3Mc0TVsYSI6HNT9WxIsz6GtHMnUUjvs9YCFMz0dGj6mzq/wu8MBSBuks13QqQmTM+aBjxr
90vF4CL7wQZIszAkS06r2SKkJa/JMjJt4nFLgbgBl1jai3SkftbfFGuh3fVcVwCk8+OJQmLfKZao
AJSacW06Rens5n6AFW8EWzPRmJiNPZoxqw4ihintfnw/6fsxt9Rw2S2naXyR+RSvUP6IgzjI4GKO
NDHeEcsOrw2ju4hvIxTjsls2yUq2ZgrdlGP6ppTMpQQj2C39DYuwOIMpEj3+gAS4n8SyCnCTZSQa
5LZ0Xc6J5xkkAh2lVDsRYst5c5YDSp7IzRFK8VcqKA/7x2jW+aYNNbCzs1bLrmhnpXUJ9y0RHojO
D4WmqBAsUSWnRpuMxDLibaQGuoyJoGm4L/BHML3HkZIub+M2YPRivwawrfDSxHjitx1UNUhLDaf7
1unNWzzoWNTIOxWEWWc+mglbohieNBVV9X3vNjH9hBGya6IWV7a51AbETnOI3F2zVqIwEdQ+Y6hn
wY781u+LiOYHbrJkRgT9m7mF9Xh/+bD4y0ngr8ou+j3RYCqoI5TgTlWvbJ/wkOUbKqU91jkX+Bpc
dow4YGG1WgXS2D+BNDOphhN2KLtT3GqGS1TP0ow7i30It/ddUbzTNXd4XiUDjGEBYmU0ohBaJucc
ISqiG+SQmfbRGG4U+Y3dnRqi+wNNz1t/bxNwh0sQRFgF1rjnd/BVhGsjA8o1XMi7sRNS/0c+x+o6
wcbYJwnLYzXQqkhc997Tx/idWG+zujfL6VhoxG8bdYYec4F+ByEznoZodaHG4bFb/Sqh5ESA3WsD
DUB7gV8kJkP5rSNs3WDzlNmDONW+4vX15lMG0fLgiogCvf9H/pVGjKtDRAk7oPneCGzwhXy9U30W
7yEfONBKT3DL0jyaTniSIHc7nfCRwp/NYVpHJ0mZ6cWlAVMdpNSN9HK3B6VCmyptmNBDnhVkk5GO
371KLEZZDGMIOUAL6r0qOzuk2QJYyd1eWapYUuUvQMlS5WwWbOcyQGH6zcQB5jKPiyFK/QwyFrxj
TPnh5nd44LnuiBzUsUQ1q73XgOVK5Ln9WVTxWgWtGhmc3o6fSPTSXvKDwLQUlPdnxU8yHVPAMG+R
RUKPRYuSthiAebTi8aWxVEYEiJLtuL6v/guui+iEH3QhUfqBFZ/2WvezdFHAuG9+XaMf9YVzNJDm
LlJuDmrCPdusnZFfprSBlGBZWGDqgpmoKR5Co6m+8vAip8NracCpgLKlpYGbIY3aupW2I/J2lKCP
/gUCpsFL2ORHlYYYBsaXTrFQyiPTn4XZxwBorVRHfeceWp0o4BdOUxhFElCwg164NpbYZUMNqVaW
JdCsXCmGrcOw5JULeS4R+owd6oHe+L0mu0ukSAVM50MD4GAktgnKO1vH8nI7Ksf61LwRYtGU6xmR
f9Hz7iUZ2x31OWJ2f/S6gm3LVYAtr7iN+7ezJlrmWndyJ6+y8xjTiZu7bTr7k9pLfnFynW3+nise
KrRvj9WtpevDAGsy2m5FzeaTP/G45P5gzKt6cbXc94KKCHCW/yTt4SPWJ4VyZsf66kunRkU6yj6k
DW0XEqroaRDXpCieo7HGhzfqSfPiLtabu3TS8el3TmfS5Usyv0i8ualbTtItnJP0UDUKzGR56Lp8
ckh1PpiUVpzjgsFLyzqw+Gck8FdlUfvrOm9QDde061LKOn6KZHpyXA8Kh0cVILBNYDQb/wTWbdnM
WE0s1SxBfvvKcFcNm6Mf+3LzHh1Kfk6d3RoSVd85WDQQC2YTjfq6DL/35/oS0rE5miDS/Z8ezDIK
stV0bdJj35UUiaW5LzpycH492Mr68tS/Lg6PGaQ8UEpapQei5vSpFl0XRp3E8FllC22jj/r3aMwM
2rnFEXlXw+xCwXbfO+DsSaffA3WrOvjiOCz52YgkLWmQ86F3+4izJ/JPMTUS2ztpHRwM9+TOwMbq
U23TXDpjDZR1FIG86nu4Wdr25XLp7iia54ZNQb8FW1afzZk1eBPFCJvrU0uYhDQSS0CEIp9L4YKX
1DjFl763P6ZAffjJdQxxQZzc9zuhVqXiSgfXgXjuOldNNcP4U/l7KBrVvbhwxAhXM79otZDvmloP
tq1/8qg+pScoKdzRPwnBUUAymhF0jcuDg1vQGQwgKaG2C8LuOIacY4A+ddjoZA44Na8Iwen8LyDq
gJOE5WMnGbKIFPv4Ji8xpeX7HYkbV1Tr38zOVrq9mC7fTK7wyUamEtO9vl2/rEfk+AtKeDTj3pnX
zFIQRSFOfupkfHSgRJ9p/MrzzB/A1+QrkGIXy/zctPMrj6H81kIFK2NBemMDQPYwv6x1Bey5uZWe
8SncrL0zvuArRr/d9waxnmybdPG7oLq/QIui95grXPJsWCgrtm0iuBqt0Fd+tIhovR9EFp83dF7X
OvIahAyXo87cvxxTJXe1ZyWPADFjylI146JM8tdpNmre/mLSXoe73Yaxu2baE/uAvHFVExnbZO5l
/wWZBKeHDA/AkCkwE9gi6qL1/ZVS8Fuv4tPsWkIS0hahEi0fIUTA9UB0cs9Fy/om1yz1fqnaBVoc
ZuZjTTvIqWTCaS4XFbzXWGoQLQehvfrmPqbhFDLygJiTx2Edl3zOSxUBp09fk96tRZ0xb9tBo/1a
6wB1C7CoszRhrSFOjhG0jj0SFfFCZLCYx6EW7ddqSp6+VP3E8j0hRqMxK4kEtanCpwvLpt71hc66
86Hnn7HgqUHyzkIiLOQTv3fDmrGbW6PZqjHFU23R4bIngVqlse01/fYr/siis/vpfdT0mtzMt9UE
kA+ewJqkjGyDCUpui7DqlQRf6Jgu+r1aUPnKZvNtEIUs56PYSusUvZShqtqx2LTQlNeTB/P8ELAl
SicCs32Gcsw/g+CfccNt4EpSXWLIpstsbZ/WwVAM8eisttdWllIeIyYTh4R8oTwWGJE3E0jYlHBb
mTViT02aBqcg7qkT/hbbvs7cfEy3JKkjpWr/9yuS7uy8nzlO1KclewoUPksEMGtzIWSWRLroLViv
8xk3uBxZgT/lFRoMSBA86vUIz4Fv+r/mubH44VDd0BH+O36ZSliyGSSGJsiex/us4kNCetLFM2fp
H60xJQlsQGJ1yyPQcUsLoU3qBvb5QjhqNznaG5AgDpQxO6fBXASqo4oEXfK+jg09tZ4v3MHIYIIv
Jvx2ViWRA9DLRpBx41F1BWCQQ2ZXmc+GgEZQwWlSrlr+tbvbNbbymcwuVar83/mpzAbgUQubyce7
luF6/THYVVJebXDWOj5BiFmcVOYVVCI5R5E2o0EfN9qj0p8m99LBVtLCofW760oadjDfyGQGLQCg
PF0z751xIrLiBUg83xDR4vO8d9Ag10aKsP+wMhRJ8B5JfKv/E/WX4VL0TMYUYoE/3RyKkpCLL29v
uRwGBh4hdlk1Q1Ncgr0/LoBdMotpNOaLxjceank2YLsttVRrgcgj+sBHTCNQnx2uFscyeKlt4rR6
1bif5eN8mYdWQdsCVNZ5FKPqIapcaWnADu9EGMG3+0S77Z+11TNW8DtwxaWWAnTKnWVBJ9sRlD2w
FnnfdCABaxeQi9PhkOTWqDDkDKL377/xFwLVlEJ8Fkiq7OtSGfUYbKQwSJBvdVmwo1sqitLYkK3A
gFGo4UtlEahJd8FQ5pwgRTf5t+7DMf2IzN8fPqL0sBeGsfwf2R+JKEMqpDIy30iXNp/Iy8vCVeH/
N+nMDRr6N8g3OqiOBUY/UbHIVdFGf0B/9v4dvNC25UyYP6MzVoVzsFwV5B74M/vzaSrpYI+YWDw8
byKTvXH7W/r5gn90JqxaZsHhAC5TIKeBe3hpk0TPN9rsjFx9cg9k4csK2+5CdZsvDnzuY1KJpcQw
1UkxKtyxtLq5V2YLEQ6vK4mzBUcovhvERx8x8/G4zn08+ZTkQY+vepuKXpaBEJ8AgcOw+kFDRuFT
PGiupit75aX5FbXCLwCMOZ8ejXmtLoKNUB+SLq8gaSCgIt/snwCaxC6GviG/vrOY5hUKP4XbNXHI
UghOu0CGq5a2shCwyK/qj7u5oHsuQLgWtOrF8Fi460T2i1F1WHvyPvfJWZBQoAId/jrykB83ix//
+6M2t7SeXRO1ZRDexV8QymfCoudnV8ailL/3CKt3Wu0V2cvDkF4IMI4yZW8p2eGmCSK9e0lLBqI9
KT0hgZ4C5B13s6sFJX0QIkemNHsURvS+otKyGujpB+xPZqBnP9Ju7aie5flUYKqbj6hCWe8Kb6Hn
ojsytMF+agsS4BJ5ITBxgGgTws27usgKRtyQP8j8XoDOk+nGgOf1LWsposMQQTc1PjGHNJCg0I5C
oKj1kEDxS6h+10NSGpD8LHiEimqXRQckZJncz44IhtLIIMd8Q+jgdY/jAyHh2mpKbOS/Wfb6x5w7
uoj8y6LmAENz5SCNT/lHySP0XUZHnZBAvBpTvmoMumIeJTUEzNmfouQ+/FmBnZO3IuqUZEulhoz/
Qhy7xxg9ceDqf0aD7fXnH2d59z/emW2iFRJMAqJ1TthJv055Q0yeAjTrWm/A4n4XcV3L3KualQne
vehAORKe+4sQFdAlFJNJnj7t8+lwjPmtT2iRrCSi34pI0F8Bu25cmAVtfv+QIu07TwAosat7ZaTD
0gfp5vE4S4uGeB9UPHfIZeT9L7Z6knmkU7Ln2NRSuBfdOtZBB275cKUGthFBRw==
`pragma protect end_protected
