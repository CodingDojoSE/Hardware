// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WU6QcJ81rWA71i4KYooraTWvGBWBtET7TXxNM4dz6+gT3WlI5ZkaoEDcVUe/MkkD
mI4qIthcHZC+Q2qusW7wefD5J7x8lJ6/oGoXaj4BM3jr/3WZI2sdBRgwWdjq+D/J
ACnnP4Tx/zRYejAW+3i9jeqOQp1AZCYkZyLZnQW88q9n6wSgDnuGDw==
//pragma protect end_key_block
//pragma protect digest_block
TwnnltWAtG84PnDyGuvjlaUqdkg=
//pragma protect end_digest_block
//pragma protect data_block
ZXi4LV6XAWCwl2mE5dkyW3uttCP/AExHYWmO/n/MbSLCjS1Eesn2E5gVn7P/Yb2Y
RmGIbnFt31SU9EdyXypInIwxpE1XCtXYMGqaDqDHADIiM0obLMmPvEAhezRbzBW1
I2pnvgebu/bGOaVXtO8bjBFzb0OR/d2CPu117TTQ2+9u99cXMuW0pliJ+97TCoZe
YbH4YOxvtU6+8HCDgkpYGRbJnxuPJND/5/i4Vzv/9vZpLLlev+apk0KRrk7elzvz
jrH3yHLu/Xr4d8oO2ONHi7gXSJlvkrjOt2Yx9MMQM4BnBRqQcwbdDBMppdBMpdAf
ww//6b1Ejsk3yLien66YdvoAEPna+Shc+F688U3qKajkTQMZc+3QQ8jzsx493nMO
meCrQtLK1pVqUP+B07kqXMJsNTMoZAFZaIp4qMVtkbo5lkbMPiClPQpDY5FwwE3y
ARkVtGi8LweU+bT6OSWYEjQBMjYwKeIQFFopGEyLD+T8fcYYWukrALwGo+2VtYUZ
d+nj4Veq3B0DQgyeSoGodXRLa5HLlDmxcaVnRdJXkHP+rFnqxWkIloh1XjDEHELz
eOznq5tHFUZlDeqDmeL+ENsGMeQTL39qrYmoR5d1ggePlnYdZOW3Ks0hu1U3U/iw
OWttM8JKwePCCXURpBo1PAGokuhm84t06ZJbK1rbrtAkskoY+OlumcSIgCXU9lOK
+ZGiqcwU4LJdl+DJ2eQi+zcWOvfw3Nol6OOUtwqWYYchWxDmVxb+hex5SwPXSLrO
cDch1ZI/he+ulZDNV5QUIy0RpIrSW6u0bKem7tbnkGpOjJiJx2XT+hOFVFHaCMSy
RLFOW374qzIcGTNUXS21LEObSIBeHsTVYLEr34kyAEO7K7ekEThkruAlOoob/h8u
1lmC88Z3L1/HgkczAahPUEK+RL2rRDikOBnPNgDnF6EENzoTrutMCcVX0NUCbz8w
wBXBFa2vVxJeBJwGIz+aaJaqPQdALvNPccvsEf2plHZHHYE//tP/KDdN1oStSKu9
5wld76VqGZKZY3zRtJD1oAcK2ngml+o4wXgJkJNpoN3AQVjDyAMIpDnnoeDzUi/8
8hQ77YXcrcU7kQkN5vlvoA9xWav0kS3waKee9HcV5XQwefErVE6lmnNstBJxECxD
JieEGsCR+vzn0s4Gh4O9igcqRA6gQbuqLQBNEwAJksDqMhob+WP85LXJDCPX2K8c
4WmuKbm9BH2L25FzUGmVcVRvX2ul8wXJ77j1CMkKKv5FF0OUwv6++7kvtfwnrghl
sX1nK1IrdFN7qxHZGAB3Y3rzTCh2uI7+ifwK78QjAhgL3d6FiLDTRLCuMNKYONeA
jAOl8JhOSo2TlQjOtT73/zBph0XEJRte2xeBJWS32SsUhQO3uAEywvXsA0SnNHTU
+etp7gDbZpMsO5aPwSi92CF2wpwcoQiS2u/STGG5Gp/en7EIpJ6G5ib8KAu0o0/B
7eo5vnGvkZHmIENyQO7Fe+hSc8GbBsDgyDzLhnQ5uF2oJTET4+5jCGSmlkEN6XJg
5WrwGYDWm4bXX7q2F4ZCunY/K1vbEHUEH/bG24bQUzh94d02aM01Jb0Rt/dqpgCL
YMXqekoks71Nckksu84iZodfnQBxEQ2ecEbizHq9bty4gxdGst3scPBnZL6Onh5J
nILy3xx5AyF6yLNM/lzEK7icohX+3H3kwmiaTk/Nmdm6Rf8aXWPJBNWTWA9UQowc
z36Z3+Bl1SvzZRzRG9RkfRlPYnWMzaCpN2PfH+5g4HneOFbi3Rhwv7p22FhA5wzv
D4v+6IvWrRJQIsUHuhlIGMFQ1z0cgnOPOf4Bu3EmiUH3XxD8HyOIdyI5mUTzRldr
eZRnuWZEgC2gaF3rnvPJ6i8bXDVq1HfluCW7dhRlNn/TSmG3bI+0TK+gQt4zrVBt
NS2OYc58qtyPjOPMAzWE+A2P08qYaLKbxXeaxHNQ6mSiZmFDkJ+infRiSuSNT/qx
QXdWytG2NWfdK/VPZymOL9ym/lVcnhXULHzKkHtA42MxfzWxqT0d368dyOvgcTBZ
aOcVs0Eg0/9hjZZSI6FvVbTsLoJ9hMmj7lEEpSC3Det5oqDWcC4IUTDMmFf4rLu2
2FTu8xqynH4COhcEoqKuqEMusC7tGHhqpI/p+3oAvCY8vH4Se0KGnt18zYb6pfBW
i1DzXAQQ3B1HbC+c7djqXn2qHqDmcMicIH5VNAA8YLEG0mXECMpGRjyDtaJxRP6Y
vfOxrq1SKMHtxVKe2auL/m0BM9fF87Qrys2XFzuunEo29lRvz8o72wgEBnThrD7O
QfyzHyVzrBCwCYKWkEU/BSx4e3pAdRv/bwxCOO/XK6J55CsGsUhqwnRZNARwaizB
kdzJgJxpH87qedWY03KiGeRm8+cjE2D5lAZ5/OnV1CI5466vk78R23ZsNmFeBBqd
f20cwTnDRnOzP3ImqdSfhkuSCawnnzrnHaPjprSERgRLQ2GyEtRj78N79AxTrMmk
CgivlVABkTW4yJMDSTYNCjAF1PDg4Zp/gYfhqps2rkkNifLIpU7hf/uXb+JaDktl
2LA5UAn1Qv1txclud6ZX3V+c6pgdFxQ7tkHrZdXTtVVH6RjwVn0BoRSMEBjs9xsQ
LtG6pr3+hI9HN9npOFE+4XW0uyt+HTrJUyQrp5NOJDS0izROTmbt1yeS6tBDucOU
N8yzZaqPTi8iYBFbRd1YqGfoBOzrE7ubS2+Qad/6tshJnkJcmY66Xl2T4jloparC
Lg7Vj6GrcwHa6oy42Me0EyhahUzDLbO7fD8yej0F3iWo4addgJ80IK9RSMp+yYca
zYOfDqia9MCAriWI+B367mWOTXsYeJZMdLzPWXp7sbUf+MBmdaoiUpx+CrZ0iNq/
nTCtCb8aCj+31lrcqIcv1kOp5I7QUz+8B2zPfuV2vr3x/FaqlvBkqY17O8mq94EY
1fd3hdqlb277aFpmK5ORIwcxVgiNfl/9xwMC0ZAJEAJ5+gvHqHCDntS2QufvSa0A
Az4DbkVqtBOANLTtBiLvZF0UKu+NbG6T3VSxu1sGJRWeCza7f9lww2SxlTH4J5eI
SGW1Uqjhacp5jLUpnRK17NFOfnY7c7kZN3rjszOHTV/OqGTf2hfa7e0QzaaCNcj+
SWAmfLG0tTDUr3W9D4gJ6uaQPBuU9ibH3Fkf2JBpxNLZlsPGKdm55yFpYRrYWNeT
heuQlov3FAV4O7Wgd487n+VxP5Xp27PnlRGxsOqKDhAjvbQiHPAZP68OVeVgEyC9
oS/gf/HmWLxJZS3eloMwdSZ/y+A5LeNyW1JPcqKGVCYiB09wpIro48iwME4BNV7d
6zqffqspAT1ikdunWuXj0BYWwTfkjGINPgEpoqlfFguH5mwdlJ9Qvnff7owMT9v1
MEqTQi0PSYj6zIMXCyCmBGUVEusWziAwlaaKVvhS3JoAmKioUF0mh6irFWAVzPGm
KwUf3H9fuPfIpiH9pY9gZFeOQbxMgAJ0Y6KfHPAIPkz+UN1gIK/KV94j5i5F3crn
br4YV796uD3UNL5+VXREdF37MteogASfYZFGmM0uSizi2+fQOBCY9lj2flRrCXmS
qkNdrm8SFLFbaWpizANNtOkzB/7fm8unKD7G53mdTKxXtPnh6CQEdS0nJyjJCUh1
GT7jBLw/4WR0u+hx3cQF5jw4FY5jPdHZErwmo08aCPRsN76woyhNsW3kzU5NnrLe
60Tptqmy+dy5yiRqFQ/1hErxtTd4jaVYHqzMH0A/btfeLwPSLSM8cchbSFJaHMHP
hiqdVIzq23tLhPTp4Y+Sht+QQksGgoFWB0jtUDBuxw8KxZGMmjxt5n3vu5CWThuD
i/TXf13rRCZfKTLf5M9sqbOSkxEYeeXoooSmov++oRw6xTmIKkxEhgKpauKSLPwA
TGD7Uy8vFjbmovzeCFAYT5Za5EOOJ9yk2nbdVV4ipv+ROUba7lhtH39CwH+sbeAM
KgOfIKDcplWI0UPV3fvQZwwbkz+ETCJkRaivPHqffHnwxwySPPwPMy81V1zg7AKk
i9onb18WfcqsBehfv2lJPzrGNhfbVEUaTTX+SQDk9Z4Fo4Dbee5pRXHYBU/a2Y+5
DthdFz1L4/zwdln+BVMf0X/XGRWIAzEum1tBbUlznwdirJgTYXRzUnq6M2ogD7mF
31MdaY0byyk720AoV3Rp7KHzRwjBwxKRnCJqX+fp1tDf+0goti0b+m+UE/Sd6DN0
HT/tiM7tByr2UIU3oz3nZgxUjz4SeWHmet+ghVoSvr1lLTMvBbansBN7RhHHCR7A
eLpQASK9ml/UaiaR583XWtsVKkhzX5WgOmcOXLNMQI87MtOq1yiRjU5bfNHXcH/P
bENdd8cFuzPJ8Gi19xZ0s+SdmsuxNUHCWbslZlqU+yDK7rmEzTLC05jDxmF/Nd6o
ig2Ake7x152ec+g/uYPmlvgskuMpB13mt0DCtzxlYuzYUxRifmLbomZnq+XKfbco
GZMw+qV/50iK1vJ46EddTS1adspszRmmsy/21uZaNoMxWxIGZ1ZUAQ+Uk10CNoEh
GvnhYxOXTy67WWNPLo/WAMwyNJ2v2ZZMWBPyKhIrvoxFXdjmkANZs9Bvhq2ws64a
RMAGQW3rkrWLUN7Y5OyvE+ZvnxdajP1Z765R4gBqXV8LNq86T0XwwzBIcH+tigOB
mdkzgYS14zOAqJz81RuK6E6AAmJn4bYGO5w75OLeT2XQ6Iit1/nyY9C5SYTdOMrW
XasQ3Z0kUrsemxo6034j22Z8NtZ/EVsUwQZLsC7Ah8T/59sNt2379OA7Xld9Cy4K
6oQviLSx+5xazBTmQVFTP94SNtfpJkD+HB+khO7oKJSB/MjhB78I7qaZkT8khhrm
k0OzfX56Qh+4r7zdDWgC1thcb5+1M8ZsXNK0ljAt4Pmsd49NoRaU3RXaihTvhcZp
sbWYCcYicLpHGMe7q3JwdO+wTDCSzIowmcClp5cyK+lDzQjUgn9gR8XJ9uIeKIz6
yYIvg9tq5XVi71P8/1ARtEGoA5pOUlRfKyFJJFM6lqOd9JfN+mRh9oR5RVtwI+Mw
EufJ90bK7s90jOpnV/Y/6OIZSUEOZ33ILAtvJtZVkomWXupy/h7+D+w0BWblYoR9
HisV3YGv5Jdiex6nOJZZRL5IUqLZNoZXhyfxbgEv2EQxX6LcR/NpvX5j8oziyxcI
X5vVrFSP2qREkXwX1zb/3gSJSoFlTwGVMCIyuZKw0jMMxX4JztCachnjDknghRn0
9oWE5J9eDP5Yk0KBHaBEH5xBh2X/ZVIYs9OUu2l78RZMo7ERd9dug0qIEMs3/An+
lDRyiPM+deS6KvnSW35aqrIO5o0cGZo5L5jqcwXUkruAKCd0X0BhWuu8+uV+bQ38
3zmdNxZotCvNVhCS5yePQkmhAZKSeQL+Q+aRE2aPvgrNJwmPJN3vAK1plKAFdFAQ
V4wq1lxtIHD42sCd5ossXyHGgW3PUZq6swIUSh+3NVUwjDtfkKgxVumUlYLZ3cqJ
iKeBFrJZn5eVc+3V/i29ECTDDTEetsWZ6lJ4aKsMB+ZgsqYUnLd86+Hrq2LMYc8b
ff2l27YX45Xn6dkComQqFtogeIeF2pm5WmG2eRv9SH0UcrHvp/lNN6Rbo0BAJFJz
NcS1pZdBUYn9SBXht/iFkHsiA33W5MmObIFNEPbjL1zNLkvq9aJQwXG7H1DnwwtS
93C5v03IILLjiNwDo37HalqdNjqE1awdPysz5dncaWDc4m7U7C3Q6+1GMUPAUY5Y
tV/39Dpq6hWDDsPyxk4ejwkl6ohRICZ7W5Njs6JrZzVbmAQESBsaWPXvuQ7fQxqj
QgyV80z8dwUjK3p1LimruiEq5m3UceOV20HP4qCDFxZFE7+i2eTWbfSAJ9txM8NC
ckcXiwidhywZ/198PaocmraKMGcNY+JsL6Va02wQKblSVyNKwJI5WrGMaw9YShdJ
tlcsVK2Nzv8xEiuC4MvxE5LlxLK8HpabrbYp6bQVRxPYDEvLGi/Kh0zynEqYGR1y
448B4scILnM9ZvTnQihI1ksRmJHawBulXuFZdAEfdmJyAGrnkylztwB6i4uL7dBI
VCHgL3Azl+AzvoDSXWQICh5ISKcBhGmkgj8hluavq95Q3wZiK4lpJet26way9KJn
AYqC1464rvZfekwVrh6TKABsdCAm8vcH+xu/7UKHW8++qaDgJTPCg3UAzhB/kBCK
DMGyLOiwUXW5yaLOI5gGn9JjtehPdNOBpPHrBaV56B6VfGsYzsf8Miz+kwUbx6W0
oT8yoHcX4jwAcUssZYHUiRVImrPqhziLpMhLbFz3cUWZHleriy1ixJ6EmTDtsCZp
T2Nb6kvlhLOmcJ9R/JXc9wthv/Dmm7LlpxVshK/UL0k/yiYGWptD7lMJorvltx2g
zWaXe8Ho45fG8KcyrmUdh4rrvyOHl3zfWoItu1yeU2n4hqsDSce1VNJILuOnqVy4
ebT/36dTpM9IHOG2euVXrmNE9w5rBTCP7U2K++yBGs80FnCWx9Hi1u6d5xBJthhC
5CSLJTYLjpscJ6+SXvJ+wj93mln8cRTOnMGCZTQTAyQXY4ow6hSCvO6fzlqmuvOl
q9kiUbuxCBs5oA+QZP0sRtTNjqzjhDbQ8sE5BpNaKIPcdGFWhQSPC33nRJaJXs3T
y34fUKamIdKu5b0nO9MiDudz+V2+9PIAgxj0kJeFh3bNd2Cw8xti5NRbiCZYM0Pc
YVeOdFXHzuvT/qpnTDaqH+SRJMTnvRq9QZRK4LuaeIUv0ts/lm0LWH0ojxppq2rZ
I/yq51J2dL6n/k9XqL75ddCwFfrMpBAHXEqoKgH2rKOQlLU773iHyRG+V5EZzYh8
8jq8WzEylxvYMhwHPVViuZgncl3Z5TcFeLppizcGGkOAAgfMj3YOJ+6tYhPS9GiZ
VRxRObylbLP28vT9BAO/2PukVT92r/ID6GiiGmCCmXByVhW8rNLWvDxypmVKDWXP
DMwTJMsU6c/goJshHvNyo49ebW3D7NKa+UwsTlH0GoM3/GpUfbm2f002foKD5OEu
ckh2HzOU31nX25Rwc9PecPyXon9lh1ltlNPxzB4xgH4k9R0wPsKc54E3AcC1Toci
oU9u1rrICTE4ILjouPppwqqONSBoRlAzOhUCZBkYbaiWbXStTki9PqxXJq24+KAG
JoH2CRBIXs113mxksrR+SeLsKgrNsnHoL0ygTpAQNHHAiQeojFUUp+CUrmVegYI0
jpEQf1dSgQ5nxJmrfoGn0Wqzl0X9zN/UyHc2BADgCl5Ctlk6frNK+rH+P3+PQWzt
Hyzo6nzf2e62yah83m4fkIQTd4xTqnDQa0OshyRyv6sMtrbtgRkrtrEs6zTY62+r
5D9gdaEE1u7bJsu1F1HAAdOuYfs6FaPNVbKKUtCQvxkuRP3RJHMfhF9xMXOc1u6D
kJXu9u4qQBo8pwelL2YlvW/RG2L2MIoxKuGP7A9F3EK5VklY7btXuicM3wPqGmmJ
MG5JqBfst1U+JAoIBp6GIHDmPFYwRBmbWWy/2AP7RpM9UpcIbJidUbnNyK2DuVyq
xWw35ObSMT3oQ7xOeJgrWFkJpQq89IU17gDCw1m21olsq96lM0aWOXVqCyCkllik
AoT6ykBh96ypGpASIaejqikYiYsb/C+0YCDJRG156IMtEc8ZqSry7AMjECX2khUZ
0QGE94Z70AKjWwdSxqjZrBzl3dWKBd0lMBwv7bFUyw44sPJK3AKb+CkS3/a4RH1M
6jSFBhGqLZ10fjHDXUt7S6v/6NML0Okz7Tegl3AmiW+XIx4YlIN3LOIrMicSA1Cz
OfTxcK4jc7wGgaAm575WMcPS7sUX0YNGN7fQYe6eeGustoTdlJpGLySh5Peu/wuz
QgoEVSZ3V+noX0gKrWpGST++5UR5GeTvZCvq8SCrQTgFvwCWhDe8KOMs/5funxQn
/PDHUAiOHCCLb3i7tgZoed0difTIh1fQcgb53JVeu54FcbQxu7cM4MJL9yJwJyNp
KjfZpN8EhL/CsIcd6dp8vtHLorCdUxzq7UwRf7xi08fw/UUUM05qf4c2jlGhsfMM
g45o51ewTJIB+T8n0vx/nIwhe4jHA7DH1FeWN69Y3EfFc0MXSmRXp150UR4LW0MG
HwZplOntRsb8kzIZLmGzLYv9OgSPYFvNNfn9LdDlzsY80QTtc3qqSX43ePY6IF/m
l9g7dSme0+ncPSrXOSxN5S/tKhbdsI2M8x1aZ/f1qFcwMICMj4ou8YZUfYAQVgS4
y4cTvHDKIE/gWAyJoWYr7SC0ogElqMPPSmBoT4tGDnf6bg4C38ykgb2bPqer95EP
ZACai9zAJ36No2wduBlrBGRqT/ynrzTnRhKOtAgX5bVffdEgy9F0xylelA2TbYt6
rrozrZwNf9EfZHCoUz1sXucVR5rmo3zq7fXczigo6LoyNkk+Lr5LzM9ye0z1HYcO
/EBffBEdUmx1jZZ9Do9ZRWLMrMenzrurgTCtW4MA7zjRmaIJzETBiLi5dsNMNonW
w82YyZMxs2dzVCJe0CSPFhj5BZRkX9tnWp/FwIZkuasqrl38VdzTgZAGcgy+t56Y
F5KuwpmskAjSaC5/QdFotxuCzerzTb+TtpqdZCslHWm1xQ56YwQGtJVF5n93/evW
JV6Z3LBIk/LD6XADRTsE6foqf/9Im5C4QQx3VZBtpVhOdxbUo0Y36ZomO1lcWnwf
gEO84WovhKoviYkoHrq7BHY55xpKHPkY3eUivchgyW1tS2VyuyYxQI7QldT9DNkC
GtAHIY/8ykgVzmS9KV2nANjMwwXMyFuUVauh3gUJO2vnj6OwBXm1/+QTK96z6Vv3
Z9iECExIGBgpjIjiAmZDsqY+0R7Sk2jxuwwG4KL1bDtaqV7nRWb6NSKJBdaepQbX
9qbDvsMIdVElWAO9dBLGlYA25h8t5iVPwtjuuMCRyAiNb7PUkYNnZUMU72rPxuxP
hFA4tTscVvZNot/oBWfRymDBl520GgqKy+uYbYovWdjgqgBi3S6EVi4sDtm2vtye
HKeYG+UM4jILttVl/npk3jCU7hTfpr4ak5UCMxQNchGjLnL6Ss2PeutbHvFkd5JN
GgtMwxP3MH00nZikesHMq+epHEdjy3p6HVPaeqsTiMQC0m2fRa3L/wSkoLuPxVx2
CkBVlL656UkZBO6yO5p6RzUajeV7Xpcp5LV0k2aAyLeSYNdOVvHhYI+T+hJs8mlL
vLTUEJ338jtxe8Y1GNV6uhSY097QDsGr9acTXEe2h1p1l1524fjZ9jCOJY8b6uT+
axwPNLMGf5VE6MC+A888XPraAqj/9agh5EW/XrDPvcsd6t6ox9heW3TXkQB3WV5i
WUweuws0aTS/p8MTGsb86zZduQ9ejLXYvE0qQTlJ/WdJyI63nUWluz4gZUOlfvVg
/bkaXutsLOdlizn4clq9bs+PZwOLxvdaCYag3y/GzDMmobqFc4CmjRQKGG3MGHpd
lcA31T8prbYLhSbWmkdQ4vCLNJdkOh0Onqke1NlqWw9Vw+INXN8sQ0ahddkoL3EJ
ArAAJNBg/BJbFVF6RToFzUAXSI9m5qD04niJlicKI68Zfjh3v2Yl1KUs/zaSM50w
LnWvv2dVTIHU4iGXtWn+jlYsstFNdcHbJPqeHm5rjSoZobb56p2I60Z36yorryuy
RCXZqciiD6Ufn1c0Eu/ruKhvG0eQMm+2yhRFCPkbKOdqamWwLfeFD7EdVhohDQXW
yG0qFV8eeuwYv3Tl1zQp1QsHQEehZyEw+UXFxjRdXH+qOPmGo5udqXx4bEqXSS4r
tg6+dfp3Z7FXXZsxzzSjVl5dfCVDL7sVaixT6gY9J1POjPTQ42LD7DK511ixHE0c
U19ntwq8AwBRKhDzU2CKt2g3b9jnSd4RMJoHSCpPzNlkPdB5dOJqrsdgCXxfNG7Q
KKH1h4bbE0KkkqdvHonBI6xidtPAQh9DWZshAgIpEzSa6M6nE49o0VMlejy+PvT4
rlz+t6QOdj3L/I5omM1AIkfwKLZVHU8RjbEZLNXVZNRGvhXLFXZce8vckafkNIak
tQb6UpHopC7d22BgjIjrOjV0FNTFvsoIwzLacspTWBbmO5xe92orrxFWZ2um0NTs
vfnDAkB45dvIWegmfsjoX3MZHztISYUFnoqRrf3RsyxIpwJXPQL38sVhul0u6OYt
C+iSNACUkRvAWdDjpAPfkHLF45CpAkZC3VI6yjll9Kg0z24itLWlf/vQrvroOgG2
77DTaFitXHNCRRy73u8auSxUdoWRdjosxuRcAhlu+nuBlArZi6AeZG/vZzjo0+fe
+5ZxDJKRIxRzKtWhoV2XSypchxs0QXbBPZfMrqik8nUrYKtx51TusbFMcxCwoHtw
UrnnwwN6Yte2qviETGWNrhin2DEcbQq2X6YuLMQXrOmvL3Bptn0WEtXuiu+UBrc2
Ye/1s0dPatXdP0EirBYtJPUCwSK0BcMtoMkNoy4VZCxQfhBpEhRh7RH89iAMif1D
koUHrkPrgHgktFo9PDmbXOTKdeMrQqJfyKh9zN4uu/11koHbT0GeqWI5TbMt3cPP
kK9c03Hvp5Ynl5PzjeEmD3ErKzBs27vdkJAcBGwJ83Aga0b23/TwUYvfM6rmm4yf
CJlZnes8y0Tvz7p5yH2rElUVCL57qa0C42Qa0MqseTC8cvk0P4aBBuANYk2/iR6l
ik969xebY+9561fZ+FQkPcfFlBfxyB8EHNFWEthLNLvRusIJzPg+Z44gaOLWBEHS
jCI26d7rV5P05YDaow62uycO6wThfJ8zUW+JHMAwMmm8mHxNsYpvZ35Bc1Zuel6S
Vz0hW8Y/AM4+OqXAiylrHm57UjBuLc9JzJ8UhZDCEWt9BB9U1P8oL+pR45Zdrkbd
HZx3Pb58VUjr2XE7+gOt1CTBTvliejZ4Yy2bRiRVYfQq+uOP1FI9wt3tYBq0C4SP
Zbo/ZoB5DyvjFDQIE8MUpKIsKjCOoRB+hCGI9/8h9mDvPKztq8E7PtTfAJQWm9Wj
zqoiHo6KpJ22dXjnXNHrmJE3h2yKFAxp0equatnhBIVr1KaaHusxnEtqEeS+6NYV
SfkFINvYOEr7/6ZnhGPXsvmfwG25+ogK3OyfQd66XU8qEJNUZgBfc7CdUxKY9bs4
ZAEKWzXZat1FP6PIk/RuyqqN2Ya7Z4QJXzFMO1Ideqf6ttmPCQmz63pG2cewg7kl
fMNmbPvTOy1Vjz56uhTLVicoR3reP+pqfE1SNMttwqmiyJBUMO7EmlBNzvoqBtbW
pkFEGC0eCs5EPayekbJciXc7/i5oYqRjVToAQT0Y8NMqc0ua4lSRhUV69bzaeZzV
R/JChA0BVJ2IMCYIZcMykZb2i05WAT/oPC/oJt/mz21ocZX9zxO4nk+GxPh9v4r7
TyFPAkgKLFeFWu56bDUPlWzQh8Flze09MaqNTx2FRjIG/5lWwnyvQ04ueH08ppK4
fzT58bpKZgCaLFrTcw02m8VxD3em6h68vGbi2eXr7l5IiyOtiOjIn0uzjB8Bm/Pj
Uh401UWPvkMTKuqfH+puQo2NrlQ48pWnTWNIfDR8F/Su4i/3iQUbLkPahCpRY92Y
QhYeONb92l+wBeF0QPdMLL+AC21s/hwkzm1yWpVBNyL7+N9ne/nIbmYC+vKFsMg5
5KuURxbZccAyyYtlsw2dkwsFVUYdord4TlP7LMpJqX129Jj4ilpt1NpMS1l9P/wU
1cmYuKhb/Yn4bPMM7wZpVeiPrhvbeo8cmYHjIQRrNzIl2sSTDm51GaEGZuXttG4U
dLHKy/lrLxZKU0onQRvQ37mCOT9WnFnOMEevk1bqci3cHE11/Qvk2u2yI7Hyzlso
C3yQgPL4RHYg+LORqRz/yjwrDUsJz+Vrk8qqiQJfCkq0r2CihkRuxPCk7f8SpPhr
caIGTW//xAJZutklsNNUsqBzs4kdFS3CojCDaBhrYKRdfADWYcir6E9gLlc1BiA7
91NnYrux8WuA6tJb4KeXt4Isn0rcUpnILU2q+PHRsDbxbPnQ8pOkW7WyQ1zxDI8H
SeEW1TF2z8SuCE2Ia+aCqDaSMX87q5nUVkRVMODyzzEueENxC4j0WqY7Rrvsg+Bs
MUZeND3ZghuRrA4eJBycaSGvXyRkNvnYbyRN+giPwn2EHYYP6prihqEhsVJym6aJ
Jp1hzu3CxrcujnPdmGw/GvNdv2LC5xidNHhmGTJhBV2RYY5EKmMcf2JDQYEzouxH
IjeGfHRGcqCJ4ruTeJQ5ZqKlIEM987wlHQTvGWyJoNnsD3Jg1iRQ0FvPTB4vrpHt
B2d50RWRLikAG3r45n66+M74RhcjxFP2tEbo9draY6IPIUx0KYy78C0sTCtoyPVB
6hMjbLvn7V/aoxX0s0+Vbx1WRjUzFrfdXDlJchv+21s9rJpzlOUybrgO3feH0dyU
tVHf9aLmBmn6E85NPT6Aln6zRVyGsVLIaaO4PtUnRVKDL0uc/tdUm2hu2HzAHPOK
mF4f1T4PQxCuI529GIur5WyDPE6+uYHod4J1dcI4RnMj/GHF0zWjHTyO7kujDsus
+dyFBMpxlKMGXjsIGtZJddn4gv6rL7hh4Xe3+D17+ksl/HtWNtmrnYhG7tbF5Z+J
ENh9kyhBKFtrZO0OpdCjecnkQKa9W8eZLH0rO5hg04h7VAYoGstyPVn7+hQA/8y5
O39oJvP6jPajK2Y9NWiZqZgJZuyaK4SUR2ma3PT/itcVJVrA2dMbuGL1ikdkztz0
gic/RerdZ5m2sfDcdf0t+dXShbbTY7hKiSdTSaEWy90C9mghjBMmyK/IlIep8ZoQ
WwhiPor9oAsvECnS35VnrJl/jHjGEfZsW0WYPgpFesMzqV+JB3ktxd77aGIEK6lb
fkbw2sWU/sAaa+B9d6yhVYkOqFDQGdp3u0c2bj4/rHWH0dtVFiBFT1zUGuKS2cgY
P9cx/psdKIdtat2xR6qHDeBWMnUy25LOVn6JFh9f1gIqZyhi8GgF+DqU70bcocQ1
StelccSYn72IOay7yjmEUIZpDMHM8esmxE7ELA65J6FAB5LUyEdTFiVMHkWH/Q+9
1cVJwtwD/p7XucDGjjsOY3ksmDZy17xWKBFP5k9MH4nrsAc5HVNwECBjMC7J2jZk
DJBG/IxTaDz79d+7YgyrZip+/UViW30hiFBEUgHQWP33qZrO6yApQm4R9Kn5cAjN
MgiPj5cxesInWhOK5CFwZE6f9p2jDME4991l74JyPWR1baiZdatXz3OBcL7XHAs0
lrmJ5FaPK+GNeXAlLW64Miy8Y6GYElHHFpPIRHjnC9BEKkLvYnoJypJGC92HFFpb
zZ3Vq+fvZpDo4WxPQgR4eHVltCpoO4R6KijepFQTH7m9VxRhWxU/MXf3X35+/EiT
boOepkZDoT2cj+oy5qildOxeWTvKMJZaUZxn73hsXxCx8G0gsTL4+ui8pQEId8Ou
sX8C+rsyQbI6+myecuNPjZhf+O2FbYSqCYv1txUl519CQBwLQ8vx2OXqDEUtWDw1
P7g8Y0LipkEKmOgHw727eQ87Q/2TF8kjTGXlYM5WhN/K0mEFoqG+WFCoETdW5J0b
usHxd5f+wjOKYN7XBytqSn8/2dJz9G/3SsUGL3NVdA7kGNQUFa4UjbX3I1xuoTVs
oEEYWj22d41eydmRMHT2DMfllZsZHA+Xls7k5SRxeP0w8DdzSTLzQwLaTjAE6NKT
NZoSRjCuMfSjIWiUqCpchyIF3MXhSLLmc7P7pNnsfK0b7hFGqvq16wzd0jpyFxgR
9FQPzhDeYZUmnsK6DSwGd7eyYfkuPuH2i0aICcC2xTTT89CCP7Jq8b8WodHcLWCY
GKUCGnrMIOkW9D5PEjYB2XM3OGjtnagquF4KoJOGR3nXtycXA3MvPdMQGHCRV7nG
QbCHoLurxLuYU/IRv3l/ZVCI5vxPz0oZcVVKrp22qiygCobg+6fF7R0yaYCF5ORD
jZB0+/BljDVEPFXLdwufTRYPfS059MQs7G5VsEAu00IRm6jMCRn49UUDsgXFcCrw
KIkGFuYsUGwLc8gxX9+Lj0fsEQjUBB5zl4LbfNjWH/gAjHLa3B62v2gjnIx/0eda
Sk4Nkh7A5i2TrsfhwhaKqevXu0bXN2wRFG0Hcz9P3SsrCwOJCOFimozIKFHCyfT3
wChuUZM8yafxZDVdLVSLvGTUKBYKhU1JrhmOmrA81t+iPFWvyZwAWwbw6559+rPy
cEh/2A7bcaREaCn4VfBRceMyw14SSaleAhTSBYVGJ1+sN1actZjFqvw2r1CJyucE
IZf2PC3MpZ6xsdoG1vnyCstKj3AXDY4Wbbu4voOCIdWW8ZCgh0pZ2Wb1DW+vm1jm
80R09F96kwURHu2AVCB4tHgxX8OPwkJrOQcMYKC7YF0HVuJ++sz9MrH0Dq8UoHHZ
Etp99nMdLHLSa1FasyQNajVLFfihQ18mE0YZ86ZSfmD7H1LEmsukwVXNcpLSzD5O
dm0IYa6GFJUvETSYQDNLlvBcy0uWxKqBuDAG614XM/omS0bEN28HJAG/qWzMQkxG
EKFp9pGfst9K2TUKxBJIKjEcmN7qekQma1CvGu6hlyozx/vWYrQ0EIlVX43EMNV0
Ighgt++kMGpFUztu1ZjAlrLg1jU/e+6MSR0757sRX7r1a61lH1/FcvkPF1WOArbL
zFVT8oJA3NyXh8yAH8kbKDnBPEHyiOvw9G2PVasNAUdiz/6sv6yT0qEpTz0m4CsH
BV1L4UrFMsoBko5Zv1yzZ7biWMgs67K9jE7NHFm8y4J08DaQ503tctxSY4O9UnEY
JFQzR2H3pmuaJ9q9NIcI3FFCSSiHtEa7CUf7A9DGlc9Wx8oxLVqFh9sHvnRdlJGU
6mh5s0DH4RvzV2CwDzVfrFQo/4fKLBnId9/Ce/Pb2hpHmpR7caDenC9mPnmEwK2e
cN/IgH06OCkTl3kkD5knB2gvDBqHi3WYJBrjCN81x4pOAoBkF4Q+bcOEJMFHobOw
G6OPYGpFCap1pl1EpP2BZQqMg2RPfFUxuTt5arDyDcMwuFQZFMjsjQ/0xCSkgS9p
x0agkRzKjtS8LX8tNBc4vD3rpsd3JgF96KEwUVzou96rzGGVsS1lNGjFtBAceomj
8xmzh5oYtPxT5rfFHx905DFw/9cV3FjqDY/o9a8y8HUsKxr6xB2U/g63CtLso/Y7
SRwIKTFXawRH+Ywf67Q2h/LOEC7HAko5UtQw9nUR3MZ5sbsMs566m+QB6MxWG2di
nkHJgCCTOS3lOmcZO48BEFLouQMbM3YIcQlac3vJMRRIz5G+O6g4aEYAlLxWhZTR
DvO1k8e4+iTzzanUtHxhKEQDHFGuMW1vdsAoknPRHzN3uEzVVTs2jO/P0q1PtsKt
oSqExUZqCWmHUcT8p1rfcmphLi4Go14eTQSccYegg6NkpQlp68L1iBJRRNcwMRtZ
5lFSYYVsjtleykX9rpdBADQoWst4h6MaepEKNhoRwhFJi+JJLy6hGfK558DVGj3v
/x8EHsJkWYfPbPS/oD8DiL7FGQoh+9soWTuUukLOD6KEIR2SvsIQR1OfcSAP7Bfk
N7n8uqtrZJQhnCUQSaWiAHLEyKCu0bibidUUoo7Z50g25cUK5mSlYLvLsOBTdXRl
AiqhRVmdFvFTTGjZNyvQNeD0nE+/71brF0Rzh5COeu/ECyJKJUpWmDZd+iL6Kmpd
C7KH+D6GA9aFeruxf+DbEZn0PNfUxQLf9qRBJcuDsq7idngOqvhCq3QGF+ziNw5o
ju7apLgDa/NMkRR67dfDk0msQlfEopfTUGuI8M2ryzb3mHdYhCilDOyUPhUZNUO1
G9riEa2DqINNmCg5sQ9+br8tAgBHk5votHG7GA+aFlC5hHdVDzeevEipQAmVvlh0
M5P9WaPPh6vSNShI0JpvJWQAlS9LxIK3BRUWaReOOjqSEJSbBhdazzygjA7/wpOh
FuTSYqO1Ngti2Orxbmpv40/OVPiNGRpzvYz14oc/njo055mIXDwcDuiSC3bE4GGD
Way51EwYPvjz8bZZI26iQ1biupzzyT8+IvzKYae8dlTqlZtzgpijf8vPnipuVal6
Z0mCWN9gFj7QD3yP+2M+I2J4KrIWPPUoQt3TAnX+GRXRxGbn9U1NmBlDTAxR4ncC
xW1zGmlQLDZumTO5+Z5qhUlCyxO/CXmOkMEPJz3p1qgBYc1JCg21G79ISYoJN2jy
gtQ9O0KJ0rnFBbBpw++6UIcBAtslmcqKjIMvbAmDGtgSQAqP+wFYJHZ1PFXmnuR4
bBYbKRv9qjXHNx68OPszXxBcLtqHjnRE4ZZ9JRidHLc1LE7Ko12/xJC8JuctLIqQ
VltEb0JvJ9sRzscP9xQsIRFEKDHzAJdsCGrOE43nbd6GOKM8xn6RKStkgmg7oJHK
+S5c3nYV59mM/rO71s0ceemnb6LUmoMYIflotAaj6XY7TbqWyBHUuYPb1Laoj0Gt
cfzw1RCarWADlyK/uhoV1Cy9uGKVOWyw4VlEO0qs7uD8e3IcepGa/8YPkNbMJu6M
W0jQxcGHWLUgTVJataL415aatbuy3G2OMmRetTHXjPEzEuMywPcIdnPF/Ujs8J4u
6+sAIMw3xz6XeTXmSlCPVFo+yIaPEtWaR2r54kuL8Qy6OCaRBp8t6n15T1/Dr3cG
PL928mZ1ddBlu5T4DXd9CpucEhbZo6gJyJBC2KCaqKLmTy/g7lUYP8UkZbw0QxvK
xORlSlZ9nFFHb5suGvCc5u1ItsBMRAsqHPm21TgWzmwXjZHD3RQ+LpWypK+Rjdnm
3JLRN4l6nuEnEokqKM69HIynQwmAIpj7K3V1GmLWTOHxm+87iFNe6udP1YHzvs00
0U/bn5I4R4srhl7BCEa6mbnFaiDXHmwTZwO6DuaPpVmUFsc5vTWx0G7R7vrVvUwK
TfhTnT+OlTQG/1ZsMFtSZ05Ro8ovN8GXlx+dux30iFafiQuJKlr5TPTPT4RobVOB
zvZ5Ew4uBQMT/aeKMw/YR253As27ij9m2MvdbB/a2bwRbD6/EqA3xZcyPCeOWPqp
uPSkpWS2kIa2ih/TLXWHJk+3AGME64cvX/YaYyA7m0OqUzOezD6Z/nBaoKKaHPKx
tMhUi9kq8LfE/5mkglpf+eQRd/NdR9an8l+txC4QGC7B2wNiyv3hzH4h4P9yzAXi
Y4rXk6c8ijdMnbhHEWFKBzKpg7CkXQ9Ns39IqxNDYdDUbcn1lJ+YEzvzRknLeLZt
JKCsfNyJRooqIDPaCu9FEke1AFQ25u6eLA1wjWxk0R+PSE0echTaoBrV0yP6Bau+
eKAzm+iMrRb4RcD5dDmmNNgpTW3pDb40WPiCAL5GGaqeQkJrAO8vqOyLofDYNk9h
sezvUJ7FYFtyG9Iz9gx/+yz1M7OPmcd5CdizQJTIpTPcDSa9JugpgTAURWFtspBq
PABkuGN1RgoG0QOebGzb6RJXXZwYe+L76IrwFAGFuizAtQE4bVvU6LQyJSJyaE8K
CMcGf3uxK9h71TfqWdvZeA5l2Z5nxxXvifcwUZrXQ0J4E2uLYZRJIFUazzB3ID3X
tCfD/Jg91wfBC4X9JNhizbzZr0VZsd+GPIneCN7iQ8JaOoH3JWJKkAJFMV/gWz7q
omWDstFrGTr5Z/4bPtOeBtjhYzXfzIhRi+8qeyVz8KvVT8/qYftNo6FS6PhRFi49
TosEouXelXOHjMl239ioL2XRYTNNCu6I+J7CF0eurrOexex9WsaX/luxn6FxU3tv
B+qdCpHRuwAC66eqUPkPOme7ymyy0fr8NM4ylIOflj9b3riDJismjHFLJ2vYiAW7
LJeh9Bi+c4Fdiv6OFkX3n1Mg94cYPmPbowZUnYJLb+5CidktSkFHP/APDjbTTwGU
0t1kZOwK8TC4LPIkbSp6bNBTvzm1d9xnv9y342QxYQMKNCGcN2YlXy8C8xwnIOvi
8fsei9EzCP1+QDpcycWvACvRxLpunsBJL62iIZRF41CxHM8fn+GVkvt+pVHzb1ys
HghmBRAl0NjPtYH7ZtJ/RBMKlwI6xZyjfheSXDAhSLOUTNp0OvP68cJXB83MyTV4
/pP7/HFUhzoZZTgH98UOHX+BvgmeKAJYfgFRGNkP0BlqWKBB/lyWLJLHmmi1Hq9t
JOkgEYachoQJ0ozDlkiFqhv59HE228Tpt0KoZFvXnn6oMozoTcTKJZVskFe7k6BH
0BnI62P3OV4eKHKxS8OIFodVbuj+APQ4tDImsWhae1+DsQSAax4NmlKXmYP9neUw
0oSxSBWAel7A/fpChhUAVydWYi8yhlK0j7YWFjQlR6UKLHHXFDiTBa0kcbwkS+re
fdOXx7+po9EovLs2Nd/UlQ2b+A9MH/N4lgPLcWCA4wD2wqGpOZ2XN112AQyz+1lU
QG1UbekkMnca49UcvOVGouqZ7Ptvs8CFa4ebY1uwZeUaB8Rg2A2G406iqSfZ6lyF
ijxuQgczJB46VBt/u68wxYZXMozRFrvQw7adVKnEs1D8G2ihQQ/KsCJ3r9h18Kx5
Lpabcs170epJKYa1yz8J0gy5gC0qVTfXY3+12MvWPgv4Txn7Gj4Cq4oLnm635lYj
qz95yPRHE+IBFehcni6IceJD1kA5+2lJIzUWdbTtJg8tsKmRlo9ZlywO7RqYGgod
xmWhq5ndJWWWQNNY7MDTR2R3aieV7+gzxR7fLaSxEhrV5/i2vkY7pAnLcrLkZux0
14GKgCwvn4ys9Fxo+5dryb8JrfEhh4eB0jqiZ/hDAyKAYJngzIREbWqnGGmsNFQq
noLfrP11xfRP2SEYO1O/KFtovX8JDw24bkDum2AVYrRyVWf/QAKJAHzh0xSJma21
K/21onDHPL2zRxCo92GFps5ZlemAEutuNTEX9Z/+0ZI+vzS27d2kwVo7A6fsaqSx
XT+a/uVhyPq7z70T1qGthtwvh42hKN+GM8SVGzwsKSpuYsG94dRV3WJSt84mSMJX
eFIGsM2jmWC8yUbCeKQqurnSyu1LyBcG0RJA6hYQ5kVk8lWvgsaWCFsAkxgmeLLE
84zu5kw5dtLt4mHznxH+azKB7cOderyv+tRLIuvX/J3aAmzg2vJU+IYQyQLADWKR
T8zs/5y5wpmhqcBLO5sIW9svPoNBijTB80B3OXqg+SI9mR+RGIpgIdpSrEII10kV
aUQ3ukYVh2vVdA9sCFm+i6r2rf+GXnn/wBl/RekQcyyU/OOdyR8RzBme6hpV09g+
qdkoiTP2hSEWdR58SR6ZDeHSMlQyWKRuVqi/YvQQpjHwVyhsUCTvclvA4y1/rDdO
KXKsvLb5/TL7bKMoSOcy5SUEGu+2hKQwtbtspMzP1WN3023rtjm2iH+jE6QW+m6Q
F01m6oaNa+WbWlF+PKJqY/Ba+20rt68xlharLUp6kYh0nbPMHwg1Ns08tm7b5OKg
s9v0Xvg60S2ETj0MiOT0B44yo0CRFDYGKv7szvh+MthxSNLApYlMM4cXKNIYF4VV
87KoFJOx2WIR2hR0Mub+7qaMRYF4KdwpGZ47FpxO7GMXVM19KZ+kUO1co77vZear
8ZxXUb/ZDPLpP/iljaMgr9dhicOVuZ2XhUyH9W1d/QdFE8IjYLvNQQyLzzBoWDi2
tlPg01PnBK7Eh4rWfe/E9B5kEForTsd5tlW2F3PPbzrdbSuHIyw0WhBGf+Of7fxp
ddhJqOU4KjR3fryzt0wCcacPdOben/cjEsviTWkeE3NNYuJnQNskyds5bSNRhfAd
KqEdlWCcQcAbni3EzHq1OPh+IaHkCnm8H3ZHe9bZ/+C+dSBAFw8+t5A8W9MlXo9X
MDHbnPxlWi1DZySUU9SLmURyy9OtDHp+POTKKSwcVsTwk3Mx75FMuNUlag1rZ2Qs
MmaT0ZndFA+Q/ZobawYhLV4rxq+swz1v0r/sAUxN5aHnMzoMmQK//AyxEzNSB1wB
NH/ls3ah1YwAmHqrm1jcZbaQhUZ6dZfceeBtfhn7ObexcytVuAzqd2F+zI/wGCJa
YnCgycJr9FIohMHUqvKNzXI5dnD5YHrc4E/sj+EmYSs7cEMKGmI97QKDB+YlVp47
lkJj6rhuKIQuW4YSZvm6L5ayPpJH+jTtFUp+kDL37YcVdFHfdcxP4jYT9i/Rq9lO
f0wU1QeyXe6uG3w1wzmWs04jUZyFeRmbXu9otrVnLLm9hZ6lSRKaG+bktcsJyTAZ
1JnINn+HujZ5ugHO+Qs+0dTE/lokrfdpWPquRF8FUTyjrjRC8liKXeA4rdoNF4rN
IeqzJ6nZi3YHZrjfG5RKS6nzvTj2o8T7tmUBZ4YcBWnlcP7ycP+5O4Sro9bDO5so
L9oexfCjjsTCXGC81NQnGoMeR4SLI9az6c8rvH3XjHLkNjj79XKWkzSk+Mjgpavu
HqPviXH0FnToadq/ZOOOmtUAHISsvOuEAZbXYASVo75EF68ZlEIaJGerhMAzoMyV
UVTbaKELCSHKCSxsF7/hte7WZFGqmmGqP4K4e3+24wXh92QbVJVp40KMTq+8Xio8
+H/GXSXtbiLdKLn65Hl9Lf8UffLQANjT5JGyFw3dF2a97Kq7+6eTf5m7h50trBjg
tPadj12BNMFdampZunbgN8S0cPWcAMB2w/ZInugSjYm3pZe3vIeDW3reqYAXldO2
8mYPpvPvCeSqK4anTNJULwaTDBbgfCEm7QGLEqNejs/nK6DxpnSrST1UBlYyuy6J
G2H6Gsrgr9AUEjkaStBQTv9JH/x6+mGSYaojecViY6l/sZ3Glh5aw2eSoRapk6NZ
gpgdnsXBBrwRpaVuaH5WWf6Q0MxLoRUmckXo5W/TNmbl0yuHrex1scIi5e4awfyO
HpPfsLOM0Lp6bPYIcsvN2bI0f8t6lrMEOVk6HyjpZqtOdhLmArXvRg4zn31te4L/
2JCm9tYzPEMClcQcAxfuotSiqpZLN1yJac0or+9zZdaIpgVkBICBpANAxrHH78lf
Fo/NQuawi7MLDOOfdkqBT4+86lqey78g7WFbsoLCSRQEraLLN79RAzoVb8WT/oKb
ijFJ7E3cObYL7hmDy5lXksmEe/pkkjA6hifv0WjJ8gy3kgAlg8JeH3BSe2BvsZRy
sqFGER08j7aX6QkYHinzBC0jDv9S4QpaqJZuSS7HhpKR65QGJVTPhJm2/rc2t124
tb/zYswWsyQFE3U61SjDUroswKImijlu633g0jbouriMM4WUwZI9zyuSBpd1xFDF
hXavWHXTRMXshe52dROHG2+dXgnFvYPwj+y5SHHqpw/9qtJb1DZx5fSz+9+nFC1i
JUJQRIJmmWUAD+cMzkTq9a49fCmaatUAduhhMrA9uHmTPuRCdlwnLE/e/eH83Zcv
U02r0Tk7HORJatujdgSvOLq4Lrq1/lMlmWuk4HM29/qidh5cGh5iEVfhRdmxIdIr
A34t0mvYnE3TwzKCmg2XKCGGkXfzB9qUOx1IkkJfYYbzl+o8dgCr8HJolWES/+FB
e+zJ3PND2Uh6WvjElc4X0BwAz9DwfEKc00x2FAa1XpTIef63mL9luFFGzTa96iJZ
uObP8SO/QshrCW34vubyvoXBEzyJcq2q3NH6HrPr18ctESVNKOVIJqyP5lm17/e4
O1Crf8Xc9S4oR7/1WZ1Urk1jPp4lQ0Q0YVTvyRuKuJXe84iTNsjcCMH4J732HwWe
n9GfLW/XAWM4nr3oWnqEKPW56uqxNnI0p1w9M8gNIFEYGOmcdzQA0KxfbIuxaDSj
ixUSe3EcAN25MPOLe7dXu6juHuJ1YYRRY/YunJ8AVgjsfZVRTpCqS1Y4T4o7Zw6f
T9sNLanlkbMV7OZJPaVfsFnZnLAgQg8v/ju9koFhhzaBQVcPRSIKv2SYNT0E6FMW
gUBNSlpZ8JgN0uAyKid9iBjexNyYKo9tmengzenPcznBB7MqB1d3NmMX/aFFTqz9
Lz9VSz4X3HCHaU3+P+IJaB5ukWIugKGsPj/EZsECjZspvgKsVYs6nl5nnedqg6TI
OSTuwtVuIwl19enMnarqOhTvWx4Ef4tbidlmz2GLBe8hVR2KsE3gshhffJi+118Z
gTeexSJk69t7vjfw8+FBInLpUYiirxvWAZzs/W3/RH9b22SHVzGmbShZo+hFPTKP
dnWRbInM1t+Urno0+oxPfUv0bZgvGM5x/kIyf5MaigqKtd2ZbgBcSstnBuHEzIa1
QfL0P7vnyaDCXKOqN/8TEU57Lkhml2EFC86TfUXj7wg2Pd7rB4sI43m994RGi+mO
1ZIOBAetbZtUlf81gR+wczaSFoU+zBjO4YyJQ828NX+coVqziFFnD4QeW56kimtW
TqNu/cOwDpRz0kZygPAUYsJ5dUWksEaEr2g7KQfDdAIf4Jbi6JCqoQ7+X3ZAe5Zy
pviaSTHjViMBKE+ENGFQ1rfJQRhRb0Mq8Rz+SuLxNT9SVDVeym3IYtfVeCJG2oba
OnydhjyhlbXbnf6quCufvYFnRDO+QLTc4YjJGZ/y6AAClx2NftUoIuWBiZJxZ88i
6JE+CsUXO69iwezFFC3+oUK9kJiesRORy5m5iRbSOBmvOnm74e0QlZwxomjNl1DO
6cEl3LXDCscWIp++gJQ8cTCGZemVjJvgAVRodU8pj0PefgHIS9Xq73Y5m/GiKJ2X
XbMcScvLiSnQfzfUsfGx7voWz0uXzt9WYIhvjUi9cWoz5/BhIhOaXirGHCZIrPHa
m+UZkaX+Ie7u9C+GhEkR8XvJNtWNBFfIWU1uYIYR1/ew+p90HAT6Ws47c2RnrQai
p5An4OVbIZaDPDeeFFkRRb98k58KlBZwhV101NfnC+t0f8+YKIfULt0JtVZsyz0G
735rFvGELFY55UbtJrLdjjC1jBOIdHHdS13HiRsJC5w+sWNZURBgPYR29ucOZOZk
jgUmOn8dfM9fPQTNQTkCoxA3/Q75pxQ/v34gjuzSvVUiH25Q+vpRApvou9m6BQpu
Nh9K+Q2lRaRdQdm/7CyE1a8Z5zZL9LqVmQ9lkKDL1mDhnVTUvk75dQU0glD02oKY
/BLfpP3U6KfgNcJGwdR7Y6+geouAIwzEJfDwOS2LJuTR3zTneUpfkXQwJzROaLkZ
xNs8Wo7J7L5fthIO36+xIb25P+6lVqXPlFG3NCIIoNNEQkEfnhVHOL2w7LjDgY3G
aZdl1gOTAmYbZ6xQ2bn9cObY30exLViUwxW8hpfZj+qRJPQfHjH6bvDEVq/WNl8A
XjHeoHFfnc92kWEHv2jkKr1I/ZGGRgVuEuIyMsZUJp+pkICW5oX4uOdFVelYIBaH
RfCIzRAI5ZUCLmOkiiLOOTJi40B+EmYQsacAmGDm6g4o1AQZE/i9GhyTAyU+u9PD
1PrRRRS77TZzf/p3lpTbV5M8b3MhyfX9EYQXyfmpDz7ZwjcJMnpeOtCIjEbfqDog
oyew+Ht3S/7Xkp6UfE8u+XfoDZwEMD2qdqcmixsFw6T8Jd6UXknDiN9LSQoX7Ulo
fWnBQGCWiJdZlTTGNzJ6mn4nKc9JBML6lZ3yfwu4wkDtJo1Y5AYBY0q2SLVmLCZ6
H+YGQObu00yjd28oxM3oHVuf5LsUexmASYJARQkFraOitCXhbINkNkpfZmGw2Y6W
2jbDT4o74v2tQSGtRGH7pClAP12woeJUeZSkw9lmCuVzImjH17mFAr2F5cYA7Mo5
/W7DFyqUbDuLz/wQS9wXajqtLPBSIWMKYytPx9uujf75+4YhiTEoAfD88MZ37aNb
6DBhXd0LSxu1HHtpQS7+LG1zdfLX07w5zp3iYaHKFCikGFIDg3b1zSOfcNhtZ8gp
42M9pDWPs0O2uOeaxM3VtP2oa+qNcejOELv1qEVCvCKNKgM4x9be9QUlMA1IczHv
ue2BP0BVFGa71CXDTr7rZmIgqO/F7JHhFlVynj8KNRKo3VuZpFjGuqCOobMRLivM
RsiQerVbe+kRCuv4a5/aObVxxIGcn4tBW0xkFgZCf8gadN8bsp2T+AE3cm/5gw2T
dLmvkTTHSpzzJ4XllaNxkoisMNX2DXX/F/Rus5PyY0i4SlkgwDqmOPaUxM2HlpPY
VsPTyBXv011DrQsSklBvly0eF/A5dD771p6WlI++DHaXOca7BFKRv9C58E6ezyO3
SARrAb4YsKBR72KVuuCt5Eh0ihYM23fpN2gCCX4/cmNbp5rpg78ROM7+5NTNv1Eo
KBrPBcdeyaR1UJIwzeQgtIWGzIlI/hdDkzvQlqIE/RXnSffok7cGmK0TQOIQikZy
Fo09u2IlZ6EkLZOKskeJMfFRk9lOQ845NQO5Sv5IuZ760qGAwoyX0ax7ydn0dVOC
OzbFNwTHkjWuzP7t7RRPZu6NI2exrpJVEg+02hMhKuZxNAfdmaAk9JQdYzTnPFpo
8s01vcsv5NDqbrpmi2fxygUxJzXO75YgQ3VlFGNsNLO+OS3Drbhtdkwy8X48AzQ6
z1rYM6q0r/FxwI9HHKxJhnHXJqsGwsVNYVpyqgaV/jdbo7dgGPJ7IWkCc5UHNfCz
5crUAkWQuPnSMZ+gbjZE8HYchi0g3aVMrK1ErI9iaSVIgksPnwZ/x1IL8fgUiVZr
4dm/7Z3NwmcGFCW3XJBODQUwRPeqtwQAhXZTbKaSm7o7BDG5YvZCvwvlTNsavR0q
m7bpwsNi/JqvHuuWQpx37Hncr9s4Wa/wBUKyij5etp6FU6p7+h2JgiOeY1pEU5ra
/c1gyiBurZFZ57p1dRRNYh5vr4TYjbOarmMZTrZpGFzjYw58hy5Gr1rA9cdoZYGH
nWlFEeU7yeCzwo12CVVT1stVVq7anGaSgnsxcQRosVHNe3GVJl6LDnU2fjeuHPU9
3qys1vEjiBmAUUmY5ZUZZbHtdK6CNj8F5foepafTn5TuOdcIuFL45BCeQ6doIHqb
RbiGqcfLfl+tZCcs+TOv6VGU1RPSi3elcRHFQjJVf/VYOhGQi+pxbCfupY2nrIAZ
65ack2aamobZ37RN96BCDjgxUKcogbMQEE5l68nfFOxbSX4MdJYl2WFgnH2fpx1/
Lcc6G6t3JTYxSWyiFtIj0/AhsGqsQBLfv5f5+HhaA9cS9fGjHMGv9NffsrK9XV9H
wyGALQ6avCwi+/sFxjA9h88T/UYR7Op8CKRdFUcyHh+oWvt4QYdtk9aJCG+G+/jG
PGoBRueNcZQKbsbqER12e/T8bVQ6JqQQTvWJrrCp2229u7gn0O7Y7zAcQG6axb1X
dUX3R4VI0EykWcsK3VnhtMgt8R3Yf7LAIxBo6uiOo+roqcxmPda4NIZ6sCQQkPCV
BrKGCnizB8SbF2yjaNBPpvcr2V9sGnFZFUyZKPXSIQ8fiSdNKhN0VMRSGoRdPRjB
BoVTDvgS1d1IjmPET/9fG1w//YTjYTAH1MaNjTkQLQ9I//W+70XSyPGDzNuaagx1
kwbn1OKgtX8jFRgGyh9bpuCjhFRGDBypIRiVCCD75yja1rj0T+zdkdMyZ7Yf4gat
bWFkDYkr5qSFJSF09kb9U7TRhRrbH4dZLVM7XBNJ4Ni4ztb4vOnhMhiZDVQ3o8Nx
GndfnbLZdqnxDc1bgoSkoeFQ+G48IaARjerquWVkh+wyibbM1vBxlm69QiJ4gc3w
47cbLdm89FG7qyOFHvWToi/BTG1LJvF6/Wkp15kwUsJsl/ro/SA5kqi2Qcc4sFuv
ZonYUs27+I6wKzGjYV7p7shVPkLR0iMEpd7ZSCEUMA5rcs5t3+QB7fLJj8RG+pKD
/2CvR5sDsYL6aPf8AqTt0abFmNfvdnGwm6wQLIyC6+LSIJNGx+Sihc6qooSGiLX4
GC+T9XnenLiKxDDI6gFxj4o2kiIhkqQh1CxVntTRHsTXnHEvF4wzgn0ug1KUljLk
+Df/f1OsMxlT6/wo0o6Zg0R0Vg03zQ0zOxr7ecjNhbQB6AzOw1FLGqnbzYHeNscd
ywAwvcIUkWlZ6+TzL/JLVPdd1g+hTJzHDGwS5HHRXI2wMQbdO6Xqzzpr0so5+uvx
+sOlHxGaiC0ykDrDyVlzW49i1uSizpar3bXL7SBR4hnGrFD15WVUkScbq8YwWqoP
bC/V3CrbSSOVHojJJKPe8c2NhT0BijsvdmKQSkKz/CpBHRks0l1D9PihmIiHxVC7
A92ZnMXJ8bJNv93Xh/FWEYG5s5dagTbBmhMvfgvtLvhaYiL1jMmKe562shgZhMur
UE7dNgDGqrnfrYAxHAdkK6/n2oIWApywvR5p0nW/ilTPK5SYKWwhzuAqxRl3E4g9
8jGRAd2FBl5t8TVrw1+ZH+F/roH5q5ud8PvzaTGzksY3N3NtUTLGMKsM9wg9/B5k
RQZM+3U8rJk+slODv2IKlgbGN7Dt0n3QfOIOpi6eaGy6UI4+dJHI7pgQ7tZqNw8B
nmsvjQ22ds5jS6jb7pWHk6xcBA2eZioV1TMn1g+dCSw7Q6+NewDpPzfBpHpW8szG
Q19QwN7QPB98s5nontHt8jrfqCviHnUyeCWnxlFA851wWvDcYMWlm34mU4Dv8/s3
hrnO93n0xHuBiD1pbD3jRQkZRq9dJM49IfSnvmx5LF0xwaJNOzczCLurLvA5VE2V
Sh+dC6QzYnb5HV3NvRmADVKCf/DRBUqe2Ivuy9dmZaUPjgZxalx1mCHCROMfnWSx
EleKPR3TrDp1uBOs7aTgY2shGQUHhTn19aADS9pW1HwhPIoaK6Sqmwr57ezKnkly
bwR3v2ZtCsJ1ttz0ZJ9VwKqKzBHhQOhld22zbcaJq8KCM58I8oPKcP3Q5jFjR2jK
lLG8zw/ceUy7G2GyPcefKkn+gtKo/pShrjRrSRc0aXyyGkhzm1+gO7UchlW/VyCk
2/su7nRqodqCwyuqOtNbz6WVoy3kGF8PqtErsTCaUEYqeI4f+t7J+GdgRwDSOtgy
p5lC2u63SMHpX8ZvAo6kxotizJTwwb8cEOHSSMhrC3VVq/Ee+Jpr1caotkP1Mszv
sWNtENI44T9weqle/Pt8H8NjjqAtbx8yPNAZ+1Baz0cYPUF4U/Ad+jWlUqJWJOCh
kEwNoGp6V7KgO4cPOXJno6WaPuVHcWOo2qHedsD2lVRYaB4VPCOWBcgoVx35nFAs
rAIOiHxhyrM3yRfl6vgw+BAlccBC80nW8EFRa76YcCPdxQgvYTixUkbwOOONuljg
2eL1KgM7Id+KaprWFCB9ZBw9lcKqOiP0Zl/qy7DMXDGB7bzlkjVLxIYy2+ivF0Te
zuSih4apoF/D2HLsHbCirS4DLeVF0ayHTtCfrwVC5V8w/+pr4e2mCsYsCAMieSxy
YBhkEjVs2WR/58jSj56IiFBj0OhTgyK2KFbigAhC5O4UA3T47xRCdpFGc8zexZUj
CzpThhmdr32QdpsIOvn0mhtiMnrNoCtLOhBwkXLThlOBT++m1Qo0ituJ10R0WA3S
F49KZv0/4/fImIVyzQu+gDbvK8Ag/YuQjJI9rp4123kgMhKFjedJXCMV79q8RBxd
3Z2m3Fnw8KvAgDqM0G909Si/d7LfC3gyp/rCvPNurhMcyi5PRHc5reK6dO6P4NRF
Ajlvk711KdgO+kxCAuf0cxANEVKFFya+dPP+KiUOZbzkuhGPF3dQbMSdUYkMSi3I

//pragma protect end_data_block
//pragma protect digest_block
bLCVKg1/gORIy7Qi4wCGFpirhy4=
//pragma protect end_digest_block
//pragma protect end_protected
