// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 10:40:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rYY62RhCJ2pSoLECNTunWMhGUws2F4PMBcvrN2spw7Cr2gzPxpz+S8k74u3rKnNN
j0664G+1YEantiGGMZZTWVX60W9hNc8bsC6phNADAt2rFERBoKBN+UY5B9mzY/va
J80Hb3Q0eC0Fhn0eLs4s199JB8typmErSmlR7bI5j6E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12512)
bS4kCK0rqG6BNz721CSdmt1s5YxsItoNd4Z5gIrFoqbn+wijnMO5+X/QTtUCVlt5
8krLY7wQShEFwSW4vXVWcUTGROC+96STOomSw1MyMNgwe/UiExCxmIjQPtUbqAG+
+Xom7N8BRkXKvKOA5N7aRxEMOAwE0KLyQpfhuF9O+0yelH63VMNSw5VPc1uJWJyT
aKdZ9RRknWSNP4VMHYrWQuefzPIA/jqu8J+r5fK+IHxzciJTA4ndt1REpJgsGazH
wvp6zMgRtfiG+6OgXieem87r/X7gV1MXfKvRcyi2rorpAn2nfA7OYt5bp8z4Rquh
SSBLmK26TMQ3eyP69HmJ3jbYpi7LUGzmHW8kJQHiR6smqI1dPf5KpwwG8j5VBZd5
tfPVtWVsYh9gfNRb/GRSZPNS7DNSwUFlO8zHXnfRnvW38FAjH+Fhnj76xSCKVQ4c
jhgrrMsitSg1ajNqgkKg1cG6oEtiTrS+epoCb1l51kBimzSkKK58K2T5Q9AxXg9B
pfOULfoKRt/5DbBGa8/MI9Sqyz/RWwXymUCZxki18zHI+SXVKJrOPXY0+jYyC37E
1bmd5gkuMrpemO0epKMfJdLAfnoG0Qu1AdvrRH9uZj/BeQ2l8TWSE1M1VjrEI6V+
gvNkZclXGKCgbOAIr778YAJXd9LLOWx86MtYe/Bkc/BywjL0eF8IviXSP7UIlk92
qeviChVBj3LNF47ow7Jzw1OvTr/lFRbpLO2vqfC/9pwxYN4UQrDT3cvGgaOAvpXG
LunK6Wna6QLEpbpxlpIlvttnAylRjelesjzLjiEgdBEX2BTEw4wNutO5jXygqPuU
+uHkKQNgcfVHPPCXfhPdA71G3kGj30rKnSzm7DYzZBr/6+c65ggBDAkAoSs0SJEG
m3pF6ZhHddoYdc9jyz2FTOzC13CGrvIDsZBbdsSdFWIWbmh74srUxho+xS1uRyIP
7VonuPE66GoqmXcgOuqpwRsD/NJbWU3YUOr+xwk+XacZFcYeVhaohq1rNKVq2xhk
6FMJ7W/kDJSmjrQC59fAmilc8zgbphQZRwx5Q4Brdp2Pxo2J0he53zysZEDpbAFM
5bMCded2blLaut0yPzVr0zhYHiZEMvs5BRjYBMyrYuRViWPN69nhRPZT4sMjXKk4
hp+P+i2yTY3vSvWnnY58CG1/f63IhdUe1yydALnhShpD57+hyFT2DPEBiyvvW3B8
Vwle+tyA6x7/TX2pEayNohmi8oClllkcQrdMxlub70fqnvt1Xu08HT8dHUbPeYG9
eBA5cIIltD6lz31iZyzykXsYDjeQwHGdzTOKI+aQEsmSACsHFn0lhZfgDkJPuzlR
wYuR9IqfkCmIQ/YxUfdZLTOHH+sm5pB8rlx2nHUxfgZbQE4pTCN91cJm+YtAqjvw
+BazqKRY/ql+2ZKJGu7j+lFI8/9bSim8Qjn/k08JKXtePSSPsNMs2A5oJYMPltof
2tVpyFQwzq/1jMxdgveJ5mJ+see6FpWjt2Fapy5O1HaTxjsy0aCcUlSBRrDjqPmI
0T3YLfqMuSitUWKLQqrn2DUIpB13hbbOHzYxcG46g4JGmdraXfAtnSane47OCqS1
GQCK0fI20MinFgNn04AKY+xoJhFNh7YUIkKGOwgScyyxFaTYnbJwnByXbZ03Vz/5
kqYZRnc/bwEFJsTyj704zpQ05DH9DQCIAT8SYYWANUtCTSajLudWvYNXt6cObnwx
xqFOkiMPyiNTiWxKbLbDrgmc+aXkFm38WcgPl1tTKOz81cbXHA/YqSeUzE9LhR7l
eSqIiEmiPoxqwHHqIt7oBSoCdIi9y2YH1bQH0vET/qvFip96hIZdpfBjhmpEOyor
7/vHxhVH7GevIQC0+Ik5WmeNXFEPprWDcR8Lj/3ven2QuNeSqBKUGJTZkr4NOGny
IwX1LZLT4MqJW5UJ6p1b7DWhyKgWkhFSLYzfo/6RmJ1u43pZI19I5cLUSaaDaPBR
fMxN4jxe03/1Abh1b5hy4yxsu3d9JzQlu2w0xQ3DGu0kyYh1IwjFvBSse2xVizpb
gJoYpQ/c+SQcSwqHV06B7OhY652Q3tmXoyZUSjbOGGxh+lRSDSGzJ4PVoL7kRxe4
149QLtbwJBXeqZWYpmbHDZGdFA/MckZS6Q4FjHQDLUSbZBHrsFrkscmoslmHjgxB
CTU3havh4vhE1rdviC0P325FMMmeLVEpNb1fonpEjh+feeNtfCLc7ceMj0TNsPDy
Mgp37XQdzun/13W8Swnj3C0uCh/LGtxxSWFX/Wnv6qDCf+rHNks//sxLgD8uE8gv
r2m5yEJ1FjKwF4+ju/5r5IZeJNCwDQaoACjEoPHUjIquGzrXMPF2E9fdfRsyd5+t
uz3Gyb9Acc3cqx85/2hlwHpfrS6bDouvMG0EHACZRBjaGjo2oSd7DfrZJ1Pyhf9l
6LmaYPD4sY8wrnXAwSB5kXD9BNp+70go3T7kilXxS+1k+SGQx+ImMiTjUw4C6pO3
8dWBai/xiIctIzC3FkUc0VlgHpXc8MG3AgkrcXuJH54lLC0oeYRcBvptS+9SkW+I
CM+KfinSgyp8joUI96dPAqFAO1I+A6p7xGjEdFteWox4vFznykx7S2oNbj5kBzp4
b7d4r8EJu+e0jFWlJcR3y86g6oyBkw1CvJzqccmGH0S5h95x5H2N1NB9R+VAeBsz
3RSweOF2aR/3gHE6uCoDIxrs83EmM0bukIn1nAvBG3Dm/MQXAUzfbQABf0H6yvSD
0+4N3Rf4DMCAtKJ2uT3SfyC/Jn819f7c3aSfKGghh4W/N2dYCWQb81vOkdkqpjyz
1EPlCEGUdC9cB1ASQcFwMpu9p4fZMvnmukHzaV/IlJnZrZCkfXAislN33GwE5X/4
/H1jM0rWtxQx46/W0XR22XPqS0429yZ0YPzKbminvBdwkhBO39pEFFBUswBDzaQj
OrIA9ewWTZVO/mXBl/QpTV/lQeHCYX/Y+bhAJMVWgF+46Ue1b0AuSo4y5Hyd0pEB
2GDJ30So4rPZhTePkmcqb/tPC24TelSbaVzJkeRAcmZr3Sf/ZAiKu5u9xCD5W1B9
Mhbuqjjsif4S7SZLUmHkCRQkQGrl3hUWrQaTqY3NKmaJ6DlKl05LhmEIpXPeLfFM
luRssl7Axw2hh3Yk02tn4mcYgpLFw2iwDWxilEMyQg3ys9ZIuxdh+2Xa8ns5QuIJ
mwYZ5yF6H36iMHfWvxf0vQ3PyvRE73Lobn32b3GQDauIQf6cbMmm1IbynYUCu7KX
nOszEyzgAEYaH1en25QPSK0lN7Ypb9mLmGmgpecV8jXbVolp07BjEsdMIE8fmOKP
+4t1zlYh+9BonodOcSQJd3Tq8sxok3JERUDnWAgr8lnenZpPEbzEK7rqx09teeMl
vxUNHCp5GwwQo8jcBnj9vD+1z5u2kwxLLT7lmGni0on2fovCAWS9Nch2dpdc7POp
b07BospY9kJ0r17DiNWTaGsjVxdjLzcDIvMu4e8T8qFe4dOrR0E5Y3DNomDpB7m+
Z5Fl1GiWzjNJJac817tthSXL0otlpMOs90I3oY81MuJa51l3pT7jDbs2yHk0Fvl1
SfBkw7T5+DRncCP5/r0XBZpkDgGJHXueFCzYbhDyKMNF8sgj5BZ6sY/mNcOSppgi
rvd/5NNyLXwFuDHRTg5LaCSBZe2ntRsjvdaOiPTn9ULeuDLPNv2LrfyCNiWvoAsH
wKvZ6okOfU0LYoJCl8qAEdTpFhH4hzvwo7BRQ05fxOJR15po5L4eb9i5+onqPbVQ
MToY865HBUj9Eqvn5fLx6itN2QUeisWsruXy8ZQYDZnR8cvkk7tfyIent11vmmeI
ZvweF6xqq1YiCWQdL920WzRQdJ1p4yMLKm4WZ5OHqrRRxUcGPG3wuAhdOyE54oeu
J9sGNNxwfUUgQqykVFAnGPSCntNAazAHLe9qw65y9akCCPZ/HlrTKwdTV2TcMCd5
EeZ1KqLnD25caAqDOAZLvbKZqgz1DSczQzho+x+hucGCIeWYia9r/k3bYwtyj0zO
zHGsjyZVAtN9rdVBNdyR1vhKVuIc3xOrgQ3AcnwOYnwBCEdQ7zmym6sHRuMH6+Ix
FM+Am9RCEM6qLCxlYsy/fFRr50tklSbmYRZeeXSWZ4mUQvclf3skmJF+5wgK9QW5
O+FrgeGEzdMKIOqtLV76gCDLZdPL3ZZAxzkQyL1BxsemRUfFgh646eXoWjHv/0qw
jaafRogFFM109LkVlI12scBUmhe5GcGets5aQwQLxLTlt/WihpIukyNcFDdzuzgE
JD9WNwRKhzUBxQ7OdWN3hKFAFNoxAXtxQbIgQD257VpU9mnQFBkDbKcOZFuPrF4B
Pq3eKIqEDXpYtvmky5VjybixEwEKCpIWOGddxdiln/Woaj3NgDAIQMPA0gGiaAib
I8L8xRO4GIvJvvJQb9YEFd7O3EvhA6yqeZfPkbu0QH6mZf4UK8NkvP+kTi+5W++M
oQtf2Eyn4BzYBiATpRxPIkMCACsbX1D7CqWoKtTt3Pea4BHddZ6GHgKwqYstcWDX
JKJgcY/15wpdJ5iMMUL3jFG1XQFFgNkaiUHT85FNhl/Ki5McbDdfuleuHPpDZ4ke
dkKQr2xB5LvBufi8a5gpGehxdJkC1CCOGENy+L+WDTgOx41ESV1NjasRkNiyi0O0
XgCcqpWMZHz9OlWv6Xl4hVDbT545TrXIYGpt8qLPZ/G4A4L7+kpAn3Sp6fxeXnjd
/K6XyzW+zgvg3+4rS4gYsniIdvDqEiECa4i1pJEuu1hWUhANmfkVQJdqOGPkVW2s
W3NihCAYeIsdblQyLlWNKu3Oold6F0EYPY89UI4AVxES6ys3AlIy0XIRw5+NW21w
iL23fjT9J04v9fFE+lmprSv8bLw7SxJy6LqgyYGlQo3Bjr0I4eNA2EC8ldMMqowr
uzoVDZ1s9DM39B9iW3l1AwFpakKiCiwRCMHTqXx6WN6AVd45ctc2Ow5aU7ErJuOd
i9haiCVsZDXCzlhXdb4A9h4xPCnVc85etLUkNR7nrM4Ch3nP9OAOjvKB9d2kVy6j
pnPKv8PdRpPSHbKpkzs/8oLtzJoh3qV/vZXwAVG1dK9/KcDcespq5Bb5HzrTLwWl
6S/U4FXgXTVeFV7qcAelRmgJrI8E13Ivq9OVfygtPnAc8r382vlNNoNg7vsc6PFs
OA3vKEPerr0upLZCDKwDxMAjG8sif510hvl+II7nVSl8rMv77nasWeein+ZHPneq
rcmLCbr9BCWnKO18cwrDaEXCXLj8p++fxNIJ04TmiX5XwK+rFzdKgRgNR+WroCtM
8lHFcVO3HJpcUvACWMsump90fZ/UBfj2AyTfPxOmQGynJcYwvJkRnGDbmiQ5nfnK
GlKTsRemQ/QAnIWE803IVUkk4h+tB2UDHn9CK7ANrI5DUCcpD9oISBxp/zSUHyIg
utK2GJHVsl42lUksii/9iTlaO280YA+5hP3VucR6KTGGlUJdpaIR8Js6bhngSGxL
HB//dfzD6tNUi5R3GtXgDTO0/AUqhhDgSIy5M6vC4peFgrrI713O5bWrhbG7MtFK
S53BGBva0yNTp0GDnHVcNj0RbuxbmBP/Ztsgn4IwrrhHQpjK+3Z05hSZkhClsLnL
0OmwXISCF5h4SdDFRQAZQjKTkgWyaZC6f0qo+acl1xORDcXZvk7Gi+qLyznTxI7m
2Fiw3XcefQxF3jlpex4Mmbebr1+M5u8u0lvKNfGeeAr5WHKJ2UgRlruJB3N25ToA
1fJ/mv/JpK58qUjeAldO/+LvXfyP9O1iDw28Fj+5dZ8Chq8mnraGmLkVDO/GD3bS
YXQ0Hl9iyMUWIB6qC5GdjOc3ZhylsSftcTzb8Ybqh1ZVlYELH8Kb++1YoQ0t5vAo
4SSZsqJ2X2KqQYN2Hn9hRrhsA7OuYMzxC3coKV6ebeFlr3EaARCuv3iBrFQ+vEiN
3PGTIxvBkEeG0MKH0VfzsC+pvjP/HVOPXlBiqvuyJsa66U2szDszsgO5WptUZEzh
L1m8we9+UBNSrcF02xWeJv6remT55S7vlZ/nJdhPuaKI2crGKtEF0v/syFfP1pDL
wa7y65rO186zvv9JlHJ5Abk6qGSrzGIs2xj2IhjiYWUzAMnKIhRT06G5LS4UjVeV
elaf47OX+mBQ+UsEMAotE+JxdesDUdJm3VaHzPRVx5li7PmseDtA+8xtjBgGfM/L
MbLx4lsMtfoAx8FuEUv5NsPHyGKXPSrwYvWnLXfKBeuh6LDvuNb0sIrMpzRwyk8O
jPGJtJ7sIGbdkpfMQLicx4xKYiV681bQvmvBDVxlYNNrDJtEBRP7tRxmPx6zkkLX
Nm/rb9NAc9m4JQBS/QTDcRnuya3uTNZqmAJobfuo1sLsxFMvrr7w8OfIGu4uix2L
zsS45ZqnzhP64b+1Vw9rUDS4q2l3vXnp6gb0wbCfsMk9IlayAHt4bkMtzoSQdOsn
2qW7BdEu76NIanocDoX+g5W6uTy1aCapam0RVDq+sTuk1gbbWvmz8XTZvo9lLE/5
Gq/9yRXvu/KSJSedal5j4Tnwvi1DPIim7ipf/C75OrSPAKSbMkP/ssa1X7BoPhjv
xRC91GS8wec9k8gBynPCRjjkXFIzkLU8wavZ3ZJod7IauYv+6/k24RdyGhYiiORq
/U1Q3KZmcTcKWQJzdEXe3wNcsHqrOKxZ0hT1w+s5yng2V/v/Zdoj4ccWoQ8jOwuu
48hLIj9dvvdHYe439Fx6XIOiEnT/pnI3J+IUltPC5hri9uBDbF6p4pD/hPaQ5+Ik
HB3KPPgDS0td0kz6/aX/EknDBlEPhEslOq7YVhGWsNVyxfdqYgRwGDESXjPLNcvv
Ab2IBY5b6ypuin/ZJHHHDGJYZwNwtjdnXkdZ2Ngpel4N9CopQ64Dy57OOPj7NDRw
ecZHwCbDRX3GgXKKlJNH3AFLMJwnrd650+ymiVRNrPU1JrjH3MPPklirgpqphfgY
cM81x4B479QnSYwP1R3i/AdJDYIETDT0nL5V26p1fk4E+q8AYICqrFziQGH6CcuM
xm+JyiR+X4SLpdux8kOAed/vOY7oqSsIwvGGFrPxzm/54SOeLJArJc8eaJn6+8Ok
W54RxrY2BmMZm20OCeduERdioJPUkwtV8Q7pjF5y8owLQhrhB7WcKKC9KE0v3kBj
3aG9iS4JdvETZvoI3c/Je6QssI7oK5NzWy7RV/QPJlXpD9DAVumMPv1i5Mr7hNL+
1c94c7XVwkEZBQZ/sHC0W0dHQOmmleFULbgKMALSaseb3QI+AnZqYNDNfZ3c8UIx
MiD4Tt2zG6MFYhR5B3kqUNrzSNbaLjDj7YxABQDUk7RANYpb1j3uCf/PYsCsTtoz
nMiKFLhcUf1tR6pt2SN5UhvSmukMGvEgzdVfBNshQ0H7yXie/Ay7hPAvlHWRywub
u5NfC+MguFAnFs8OBs4Bhamw/IQ2uYlbBisL3ZJUpiTyJcqqxlNY9vIlJJhpQvtY
xZEL00iaW4aZBtphKLuQXb0/ETG9dzuVOK5hsPU26CGBPh04q0uw1/wq6QHQ/chN
VBNDXCriF5H2L/DwAMUPRWtHNriWtLn9Cmrfg+HdR9ctd6uE6A9WgD34TOiJbDhd
5fXLHG2I5sHCeiDUbNVhT2GoPnoPOmt3M26TvJ1BEhAAM+JswfUjb9w2KMig11NY
ElgzUQPZ7MFCw9DTXtmd5BvirbjXZpp63mGpti7fTjjy79xj4Ortota0n/pfcFUJ
5zfjW14LqA0UbC/Afr5b7ISbOBrr9IdKPYsR3g7o8JkPHuTEjjN9A0eqiQS7uQhx
K0mSlFdyRMqVPqN7RuOKFfx39vVkOJe+vNdnXAWMQbtEMo1PgxTJN/zMjdXVedzA
tOCM7LxTYBNZPfzawtXwi7C0N2goZc/fx06EnSsxxWZ1XpS9VAPMfTcAzKAiYJvr
FCdm4inApYxAcnElGsYKWkvc4SWOf17l9tof41bCjJ6NRDl4DVqZBtEr1b1Amj9j
8hdBvyDThQ4T0v6+RUyAWjtKK//ozwii+BzGIvxphgjCI+YjQlySMy72Wc76hSiv
hI0ssv77uib+73yWgntzQBg3c80ayHVPCYa6CQJ4UT8fIT0M1/pMv1c1HhpFaAt6
A0qcPdOo8FeD+GiXYR62Xnp55kpNYOauuFesAtBbFgD7ynOq1QnGDD6Vm1/Plqno
WGWfYhXYgvkodb3l9APgjyt50AJYGkNibBTbEg0GLWLQY6WlTCWzZvcM6oK2SZtL
jveRwbjvMqTvEFzBAQ1JUongFnOilu9NO7ckB5iraeGrlMABJwy5TAmwh9DRHYs9
XNu3s/JoWYV848FuERxcKoF07fHursp6dmpKmh9gkwlv0j0LTeSion1aMQWvfAx+
uL3PlFBbIgEw+RUJ1cJW6ebAsAFYvqkmwpJ1TPoD+4f7Us8plHzVOaEKwj8o3ozG
ZHbmON+CZnZD4P8wffaYtkACcVG4xb2UU88r4rbL7YcbAZr89geEKdb7ZDlR2bjp
hHWD2rCnYu05pODpeMqmpt86J+d6YIgMEPGow5jJW1rPhPwMJOjTO2loTXqa8CjP
2QsuevTSQX2IummVlXAsvTWvWISBS/Q8041c0028guYb+nqz8rbCnVPM0ptfRRmW
KJLR8ouAYC+k0q22ty26jOzphzKYIlisZmBoNapvH5vIlo7cW51eedV9XMTRe/3C
moGcFlujiY33e3oonGNfJgoECfWL2MjAFLI0iwO3WCeah07DqTIJ8OgIkOh5i/Em
Z929hm/j4RY6vQ15kwVgUwP/s96nA5sBmJe3WHpMV/iR+USQMHgigG58W0rYYMoK
MXrynFRdC7Imr0znfxwvL/Ds03+tYs3hsr22N/WbBn8erjxT92zZXcU9JNzE5JD0
S12gfL19IeLEqiNn1oISLmCx03Qt6ucHs1vkHM9NPPodM+wswFHBRjGMfL2JebIT
HZW8khR7hTTnBSMOvLdolJm63OUOYBXJVOIpo4E2W0+Gfy9KAf9O5/Dt//6Nruly
3NaqKlDW5xpqmmwc3p0l4EcGNTDZebeikWwt46QbgqUAXgZqqU89n88+bXIEje4L
dWMorIlpDrksvfd3X8nXa3iB0iRHowa3DMsQSbSv8MQHuOCwA8hYLPQEPQ/8/53i
7AbPOhSDvcASPqA7lOypz2eeSDLnA4NZ4trKr6w+ZncKEP2Z+pWxtga6kZ3veTi6
gOk9dVo1sH87LDdPzfC6TjD1xV2UcqAToGcdqNp1sLYqpk4N02xchy5r6k5sT1Lr
moJ4m+a9FsP1CSuAVMFUSq1/gMAyAFYEZSoivtg2R5rVzIbRYCq84UB4BXJWRcw0
4Eyzd9iT4XZp+hUGZ3zQce1BnJYyeXFNpYHk0efLPaTe754XIj6Uf2sHLxrIn4jw
KRI80KGqScFsSq9OJm2yaROkAA7nxw7cy53OLzp556dS/CmMnruTdkpC2Sr+SaR3
pPqqWPnztu3qezJkPd0esmWiQ1g/PFSNlBFW0uy16SxnA3wdp7PnkpINXWgHm8h6
WAHi2PCqSep2M9sAnQkIveyRGl6ha+M3SKDwpdjn2x+0nsDoEszlhB7WKgOAGo1c
e/ZJ4QPHLnp2uROlSurtG3wUhCxqSG1Sfi8FmXVTSAB5pIaj3a2CmM2hTdLvlSR1
nppgBgcACGk33CbF/ZLiz2dJofaSf1nUzDdgNmR7OTZc/QWVhNm9evxrrAb4kyO2
wNVdO7l2QOsuxNzuivnNBqFB93QOExXV08D5D9aZws+BxGw0LLA1qOpSJFcDu8A7
Yb1kufGP33fNB2n1jQyCl1CgaK2093J0mo5i3lJfA7pRX2eHrYQ3PhK8TZZqi3X6
5KvZzWY4Y83m8tIn+ja8bXK6dkzwMwMfWrhvd3XdTk5xFMjasUQkrOpEDnOFeMTk
Pb3ZIgAH+hDjKti3z46jbJtJOXjFnMop83nMKFaRdxUmW1/MKVa4oIL6zOqUTG/H
apZsA6OjIvl4GeRFMjMh+g7xpYsoUU291uXqDi2lHfj6LXFXJB05uTnHLfCE/UcQ
tcUkW7NMyxyP/3Sk6QGmGNuBY/qAifjjQk2Ow+nKroJ01nmuxuiafHO78fNt5wrY
FMYL+FMJHG9/NVKnOwFVwVWZBpfRvTnXBj4nxbfWpXPafmLvgqIw4oTGoMFO0DQo
m1ED/ugM4m4axPSRHnmYt36kXCHVUgKnNMo7IUynDDTviGBn/ZLWsiLitn1zDI4M
3j05fUz+ITZPVV4p6afyCWG7NflWS6QWMGE0zVC7wYNYnZVLTiemfMaMwILhQ+78
0v0za7zDA7g0yFenDNLLeHL71BDbnMgqS7y7HgsfpJUwG8IaG5HRCar6XJLjAEfM
RYAg3+zVmUXlxo6nA4ALtTp7a6m3GELBnZW9SMTNMTtqD4oNj/HacemO1HjDnOGr
ZZ+/hhs0FjGhsO5QAmVdmaiG2ogEQ3nGpK26xWe87wM7dW5wTPyo4dovv7XnAQC4
udXyaM2ydCHuLZ+vjuSCJ+WpC4ILkPZxM4AxFZLLNeTGZhLFVXSy2qVgxRqSZYvp
J0bgeq0KfWWmd0qddDqer/q0aXYf9ojHV9CiBC2C9hxsBziJt29zXMB8HNLG4Jp3
qxJFiM1iJMc1WyIAicVYfNeUnysBW4HByjlFrq5oih0bJjnxZ2LUGP5OK/wUsLOQ
RRZ0LZD6Vek6X4qJTKwLkszmWo9RcTz4uMo+ST+C6j6OFR0wmHGw8YcCmB/7ZLzw
KpFu3em4GGhNb5xVwNJBDWSQK7fRTvozvS1OyTvKiD0Bb3ifKLOPsNa7zmE9jVqy
2dgDmGqolwmxSpmqN8sEkPJ1eKT7bNzIqjHXQNReMLkIgmUHzem1DPaP/qoKi+J4
PgMfbQ4PnVfSKPipcJcexI/0ztL8Z9uFoyAO9XKH4Z/mMxvBJyIrelG55gAhMz/X
i/ki7L5tEoRLjR7ywDaQvnSjDtIKeirCMOC8oTn4FVqJXlHmfFHzQEGCIvJhkU7P
QTqAekHeVvNv+4XaQNFDXenEHumlOcvIhAKKWdrUjE3GJHS7EdmTU5xNnN+22Imu
zvEj7jLrgj6tYcwfYr0KzYEOQ/7j1FZXkp18evwAEpXBvC45EupGc5Q34asVZ3un
FBku5hzO0KzZ8GmreCy+3PO3KIrFSU3bxMwCovZizE2CTfgnuoPqf+JQJhjpFZQl
KKYUwjfqqaLIU2RGABCMNoESK2IjtsyVukB9xNgz3rtPU42ILBi+cw39f3b9APhj
70i2OtDtH87wn7dR41vXTDc27sMeGwtAzY1KI5IRvC2SGjY5TUvxbCncodFpBNgL
7MyQaZMdvNP9w/OQkb06oHnf8R2PZNcc/6m89o3/SEhy1m1wHLgSlraSgt7F9Uh6
ryTYq8D+i6V1w9rJahagWtgBjAgUW3X5eSXgO06LcO2D2h4A2QExoQm8LhyOPPkb
UqtzKIPi3lS5TZwsRvezYI7+YJxDgw5xRlrdwCnqjNDfVUs+cIfa9A/z6bjTYDWU
PcZbPiSX7eyNzbf8C/YJFxiT2vmqDND/iZ1kqdyxexfjrqicvnSstWdZdVvhvypr
xaYuiYQNgUtr/2VePkteqEwnNnjfGAr8sToW3qIV/KgNDSy9H0vNihkTEl5g8va5
/TaDBXCAt39ZRKgHbVxDdq0WHBZ2zxWLmVkdGYyE8kpbK16nR/u6mNAQ+xd5i9LY
qsI/dEalDBQ50BRZf/A/ser+pePX9g6lBAyWoXEAMo7bqz/7ubiJbWiSJSJl//NP
5nk4bCqy5Esm6nIoJvwx5HGFkRwpbzj40cnSphz+w9knvp29o3IK/Vm5l/v82ArC
KmYq5ZbFCK/Qo5U7ve0EzN+iBjSzyF+Mjlvpq+7IfrRwRvTubhJOyIbk3nNSCtZW
olTAmNDjUPQ6B3sjl4dmNb34KYOk/ivUEXq9kLIOKy98MUxVFQGBmrD58iLR5JHH
4OT2EGU9vxKJl3e7mczwOFnsxrsOSIki2M/6KYhgWQ5lZ+yenJpFOv2+L3FdUTS8
LB7b96XjVirpJo1885+QE2E61ZtxPi2RsVRUL+m1PbZPcAEJbj84CxVEba4dkK4+
XlR0cymGbrunqtNjHha6JijBlrDY6ljjvyA+j/P4yPtfha01lWFQNTqz2AAoaL8W
FYq+7E0UHii6WRRfm3lWCZW/JjikrtbzJovKfM1Oe6xVL68rPPSvav/2E6Pgc1yU
ZeV+jEGApOUtx84bU6x+EX1bflIzHv4xxro7UAj1LPlFYoq5WeZ4V0ZOGGPBFEI4
bOZmTQLOYbDoxdD4GLwiefUEHGpVbGaTnqbpvd0I23nsc3Iilh6RsTSN6ov9TyXl
MO2PSLcp98kNhRQ7tywZxPOlnp/lljI17+EC6qmPubBO/4tz+iR/NBiA94pnvHFm
0METP/DybwWGXbfuV0wfu+B8bHDQr0FHo0jR+G7aCJ7uTRJa/Sopz0nhy/jTXJxz
YpME8JeCAdihwtTpRld84Xx/leluLg8NPRg0QqXNYGrxOM+9K6ef2zKqHaXaCT2t
pEBha//4eT9W91TNUHVB6Q2NhEjUJ12RyrevHDuoozVxsHfmz3bb3E1uIx5pH2+m
1Ci2tLj34OYs4JYHwZGXebYgcKb/LWyOseq9OJ2RtrbeIRwAGeZUzJ71TsPuI8AG
DCkwVC79itQxeuhOyk+kgnTQlbdC1fsSgVmdxzVznd1nh7CRMCetTmsZtbxoikKN
MAmodHWs2ylVNCuq3XxcuV4MyzDtvr/+DumF8EsHBL0jVGZy3nUr3zgzwGHBm8wa
fZrQUyuQ1N9ojeM1uWRZfHvaOhePD8sdEWp+FaMYzANkls3NitEGAU3x7hzQnCVG
13e+7+3C4u/Of5xKpfKg5qhzcUidSJN4SEn8VhqqvcTx6Q/LbxkS4U5Ar0L0dIpS
MacQEIRgPCesOWrGTUv6tUKfYVeZG16knlPDSwsZelc0LxsUAJre0U1/Qq5rm7yx
nEfhEy5EQFm0UytHeWQQvvW3RBK03p+5CNReUKA6685HiJkwRfZ9XOdNtABphsTn
xkIgOVYRAwa0ptkdyzmNk++BKpTPdoJ2Fot1sAw2ZmfnkZPkidCfLL0jUKHgLJaJ
hMszJA1umw4DImWRdUYcsRBcAqbmOHevO6l2fPC8b4hYyYlhL8z4mtrFYIslaHk3
pLft+U1uF4Wr8GFqezff0TWERdKEWtBOFHz/cy++XHwPU8dXlCXi6hxQ5dgQUZli
ElYrg7i/h2gbl3x1u9tphHRmDogKwmcVyIZVuFZBZbGAzFgBZFAjCz7JlcnRqU2I
WZy4s0JK1MUIiGNrhf4CYyE3iXLzhWoG956FNJ2ZsOJhHKZUzp11ifRbt3vjLRR4
zK3SZ4dGwH3Ga4tp0cskPDVXvmfzi+jlfjuuvKqf97VIjwkrKD5ORSZoCPWsHOfq
EfMsXfaW/mUojd2ZXWRB+2wjzJBEwPF/raVO26q2R/A3eRGL4X5dZjLCzb5pFsjn
9tujPJ/Lil2yWX+LXZT/JxCbVcpfE9uCiOBC/YctybvWgbKU2RtZrpuVgv9ZO9Q0
1fZVi0cXSBVb79Z3OfZ+Y7jEMscLFNQEkFI0xLtWdjlUnpgDNnjXG6LaEtsN7g1a
MXk9hkg4M2K4nHXlfkpOwnsYA8AkMRzg+A+asue5/hp/AkqSlQgkh6HJxp0PAJim
ddClkZdm/fj/YxTY8/dUSNbOJAKL+Tu+yPg0Dlmjv4X9Lhfv3HezFF8BgbSnPf+r
yOX5DRuyZUvTCeCcbVIl/k4PWaAH/k8GUV2cAIxGDaxASXmvJT00Ci6EQ1C/YXYC
g1W0SCctVJiO6639gkWPqIXztb8fcSxaB7Ib0YIH+StgpQ/LwOdLP/g8QeDswHzS
c9GXVqfht/cUX/WkMHfP/JSsc1UoI9Ov1PIzPceO5PvqYHGAAfRkKNfSV8TJ/+bD
kOBaMu0F3yU7s2FizAU4Twv3DEn5jcW/ibHyeK+/VjTHV5R8eIlhV/Hco7mGAkz3
I6dPG4z6Cvr04F3LvJSVSd3Jfg3cVRMO1j8JsRplZSyGzXmSS3MgTNPLTTEH9X39
rbKAKlwKbeQclxp5aBKFWDhYqIzhafS7cQAVolgRHvjTH91vwHDmj1SMXTuJPtMA
Xz32uLF5fbQBJJ+umv3n1pYWztCZjWfUNafThX/oe7JVmD4Z6fj9eYwF/QQ7k166
4++i+cJVnP7Nv1GOcQbqDDiyk03ExZ6pn2M/JGu6OlcacbzqzHNaahMzXY9BZyNi
kbE6n3GGpcU8oXXgIOIUIIutTT6259mUXWoax6h+t1j3B265yVYVVW3cKn0qao9k
92ABzUDm5bazO9vXy27GPJtBUmuz0qLp+fELP7KFfs6qds+9pyLSfaGfr2FjBLcG
f6wZk3s3l6P3ynBD29C4AyYvQZJiExASXa7C3CV34ZpOcpgcS3W88F9+ylmTK0h/
2USbDRzrh/u0pmvfGNNYGDDzLdgOqRgArjLGJbui0LHCgVA66ZrMmcS5U4sXuqAZ
OQEUpGyV6dZCLrL/HujWEzGTjuMGo7Vot1sIcKrZoSdKjnra/DWT795iUDGStWh9
Oky2zpGnXUM0aCE597uIzuvXwzFMKhhilAEpXT1ntyJMG72Gn7z0JHjen0ERuZ6/
j1WfKtBJF69p7TEgEGUNhCxNBiK8Fi/26gZY22jjjv9NpB+0psvYsV253RNSojDD
HNct7pcdFDvQCFCEKZqh9Uqid/0xNgqd8XRnlBQteACBfeQ/llBHxl2UdlUkmA9d
0I2GGx6m0AWJq1bOY6X8vu8Rr6Lmkpg9gmM223JAvR2OjXgflkp17EpZNvc7eOi9
sTr/BhYg8/Oc0nG/bMX+Isa/Ofo1IRHb2YvH8/AMW5Uw3XJB+gdCEozzAw2ZQng+
vdgVnwrnBhK5ySSw3O4nehwCbApTHuH1sRIq7eYYeoLBYrWGGaxJJexT9b0dG3Kn
o3naT5iv501yRlPizZEhyvgMxvHS/yfaOP4O6zfJNUDgcaEwJaBwlguNUB9u/FbM
2/Twidv/Emy/cOF0CCDlu96C6d8HehrWV4tiPU3b5XewHA1+Hnbj569EomD6bw03
1kwIMXM3GcvCvXp3d7yCcD6bfx0PKsp0gllUzEiOutFp+7Q4Pxt7U2CPjxMH9Er9
W8e/4Wx5nJoW8UdQ29tUMXok2yAWNZSLMPbLOXDO3Zw5TAfXGggO8H/EdqG0sVV/
d3CndLba+oyghXX53p2pGvULfcivCupG4mvE3nWUzogVbZQzeYdQb8RmOuYmwe1F
saRY38+oeMktBNRVRYoAquEPsHZ1NVF6e4y6QsVX2tyeF+oRd2sa3j2IeB5G6FMS
fc5ijko6AYZdA5gwVuLlRdRNhAu/cFuBloaf4SKD8OblwmZt+9MrwphOeN3IBzrR
Y7zD3IOFMcpGB5aJt+Rn7HsgZ9payY4kPpjNAHEic1xPghX1WdsalnMYuYX6L+NH
OOdVwxrLCHhJA/4UWEQSS0x2sZBA2kMEgWEavUN4Zszje5M/E8h/1VKu43flwjHz
F/HU7xuwXTH21SvgJEUE20AApArseWD3rxunMgXswFWVzTpqwoQBK/QTUvjWwYNx
HlvPVXKs6fAQO9nePlF5WP+lDq7HfNE6fWQ7s0xgTaD7mgyTVZWNIsuc0YD1GuuB
tyvhi58kmekttIY6l0bgujQ/kSBzBrVXL09sKE3bExLiuD6uEnK+ulx8QUBHWLVm
ObQvXnlN18XoaqwDloCgYqe39u0XhFlLIw+yBkrYIpmeGnUOyKnXd4dpNZptKuAX
GhuN62eiLFf6yDFFRdv2BVBuEK6KPTvAE/udVXwyRvYi0WfwrY2ieGUXhl7hwz3t
nPwRmECbsqr1dL/PjE/nP6NgxlZncTa7OKkBRAjnXMz2X5EO0LFO9uAVqg/3lIi3
nqAlOQUZ9UkyepMZPmkiHczwQUg+JikoBq4AoanvQo4sL5OMvoGlfgIo/FuYWvNx
Tn+aeZphKbcPSBd540m99uMkVbKOeZEx+sHUOMy1N/6sXUiPx9wCwRmbp3sq8uM3
MRCKT8rkWUstxnr0bFhwmDaOVbeKPs5G4zOWUvOLqv/0XfB2ynn+9yJD2LkOOyL2
6a+3tSq9BQf1oIQ5y4vFr/JAIeM9JcsQuUdRvWxX+T25+hwKm6nt3PCru4kg5g/n
ZRSuhio0MvldUvRqDssKhCj3Auf9mo+m9VWJ4qwUXbcGZt0LkP1ENknJbfDHnyQT
uoebAwOuNgPysh6bluByQw2KyxqzYlxFNxIqzrjL1xBFN4AX8AaTlNweYlqFrmew
mQGRZIr8rmzxVP43CLxONY/osT8M/jpWZvo4lSRipX+XxbjmxiJKwq1b4TMxBvsY
81akdfnTgJfm7ka725Hc3+mz/OSHx3le2PU/NzhpwLnkAgydNlcT34VYmwuptnAL
hTSkiwj3SGkG/mIA3SSrB0nNS6O646F1IHaCVzMrNXJdFoc7D/lbvWFbZaijVeXF
5hvLkhcwena4L3JPCpoXOBXhMoH5zHcR0tYk2P+Ap0GzvRAIBJLTRkx90fGPd7bs
Htj0YcZ0AEnhg6SmvF/taBbqJ0QYqVnVIGsqjcC5OhxiWpTh8WqkvsYK/WVBHWOX
ys3lgtec9x9VH1CHr5V31juBPbQ9GQydp9FZq4ODlis=
`pragma protect end_protected
