// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 10:40:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
snGvFE3jdNRjuSDr6GlGO3dmbDSI+nBIxyALD+XfxnbbVV/bLfXU+smJaLvvHOqR
8yU/umGbUauKeJrheTHHu1CW97eCfPxmenoZKqDjpj9PU5mfgcq7cFsWVUqvH6u8
QRbXxZcYTt0YS3LYeqyvWzJMIVIl5fKvI4ptB1M7T5A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20896)
5pXYHTZc2InWnREaJj7J6R7ufQ4nH39AwMuliKKjXFM7er2scq29epMUW4L0DHVZ
58k1cYn27aMOWFhKgEBr0wke575BZFuTYbg5Lf12bCA/8kZC1YnJdKQt79fWYe/8
YJ3ugCbXX/a4YvumHgiF3OGb8BsflOLnln9/ZZJTKDZocoJAGAk7DD1XUqbfmq/+
UijgD0WJ+laUHu2jvI1UwcHm6fZ26ySLlIBXW0OYIxKdnmn9Fq6fHetB2Pr00Usx
D6AdFS+ZpOlF6pRQmL/avLqBb52JtTmgnjz6wvuF/2i7uPc7yGvXYBtrNMHSh6+G
m3a1hixh7emsSQp5pfggt+uTy8RD+O8G87atmZqDryAZ+7cf6fkF+9fssdw/H7a8
FI6nCOZ7kb9OrY/7+j1yPRgZsYy3/GF5u0mewk3nnnKNK+pK8D/r7VRL4TO+Pswl
SFXjSydoUIgqs/XjtfIlGw9Uj19Utao+ucPPrLS5z6wVadiDYbEqQnYvYrWu0JM7
zTZcFmOsoAaLWRxbfZ02Y6JAzZ8FppztaTZFg+cC5vCejgYgY2VsPlN3pZzM/0OV
yJQnm+0FkDQqyqIEvqhUnWpHqnjhP44CLAHeqjZ1XycI2yZWt0GZTDeOIZL9k8Fw
x3vwiDAtczsdTtpbecrhJwmP6Gdzgri1ZDBfUzVUlXVI/bKINAbZTGwgQO7XzeIB
ulMIg0KGMWeVQuY5zFOz0uzuCoZiMuwWS+3OJoAvUBaLMvH869rDz2ZfgD4Lt2KE
SdvKEl2b0Rp32CTVfy+HgsSY9H5w5PQ0hdSbM1nNh9ZjXPAXRrexEKp9Z4zfcH3M
DbiSbpJsJ3FlNf58I6eyvI4zWxi7QtG2+JkdObhbfxfI2DBi6QD7KnTDZ1u3leIf
/0zETMQZ5AORz9LSmSVu3jzfGu8wliSKMhvB/8FGGEv3tZ7U91ogySuZqHO0NoTt
f32fCNF2AWigbS1jK7Rz2nxVWEyRYHittzzbgmfxIDLTkb1q//ilMUL9m6NoaCLW
udbdtC+DQ0jFgOa/s7oXLK6SDEIcCA6L2OZM9AwR6gcFBUSrgDwwCHZf2EGShcVm
RXavzjimzJsCyJVlxDLINLi1w3o4acsp6RIVmgqIiiLi+NrvrRw/n3BW4N4PV+qB
KdqrCtM5bXCINnl2KifIcc7yfyNs8O1NW3FArasTp6jDZlaH5nrT3C+QPl4otH4p
diT5Jdt9WDwLBGNcnD34gxj+w9/1Tv0gwZo59Nuh9LSiw1GalRxRav+4EI2kKXf4
IRN72mt6/mwgJmums7UJ3/l5uH+MQUY6Q64TOm9IpGiQwXhiznQfDEnPhlpw4qjj
pQsBzvyeb1O2mw7LzrAkk6T1anH1KhknHcsOStSMA3xiUB3NmKi8h1L9nvQHXyVN
NQfYyH/DDOJnc2MJKjmIXCO1m4ZTNv6ED3qfYJNAooBWbKRL1PNnAalmMQ2kIXAK
91LKYyJ686X7BKFJB3u8u02w7tNEMymXrBU+Vu7B4mlxatElhd9ORgrNTDtpV4hZ
S3bk2L8vaPHF16YUmR7VEQ8hFpBWmNVLXpaYYUtoRAucWOJ40NKm6HqW3ukBx3Or
LkqDR5UH1BZy9SGcXT0L/yw50hTuFNtXWG7JkIiSxMNRSmQjJZfLz+kUWQ4AjhgT
7D70vgJy2EpeodIyyk8eTmGLm/Izuv4MaIookODEyr4NK7k/s9y5stf5MHclMJcl
cCts3cOajK35mJZVlJv3eUlONEQw3EWlzvcf7mmRJSbkjFTGEc4bQRTMFAIBVh5k
Xfss/Kqf38KaSgLEWZB8QYVQi0NRmwpSx08MfnOEvViDi5GCF5T3o60uJujGmMzU
waTW3/ZXyRJtN1QfFe1g3D8TB3RZeoJS3ne5JGcf9yHk6cfK4KwB1pipjDAtjtNn
v+Zs2bYFK+g2AhmgGoP2jJIEJa3DGadespmEFDRWZ8/jaZDbKZDA9lG0YA1wkwT8
CDQR5k6HUTJogM9JHDryMEl6IOMWoZ/20IHL47wcf5LOCA1/5kvZdkmXymsvJSE9
7oY7RYHkwFK07j7RF+Z1w+CeesO5HY0FyFfR3QtAb58dmeBWJlZSfElKNy5ymmc4
rnAEMv3A5c1purJjolzVb8oq59MGOFxVJBrkNrR8PVZfk5J7+oQ6+8rxpGnOrF2r
zofYkZeg0YjjOP+TP7qcr2DodW5wVZsvT0PcRldVv3OhAsncfEX4XCdyAYVs6W+J
lZWHAZCGi2pyWaYKZ5szoOY7bK7NGj7M5ZKw07LlIF0wGT9k00CuIO7APv5v8HiZ
XNaziASUZ7iTZZBapOFwZ9zglBsKgoouj1YDZfzvrtZw+452Slg3J30rbsDxEEJw
BvcZjIeNzmPdaxmv5nnu3wvzUd9QbdCJze94WIRkkmema6vmgAtY+VL5z14kQ6NP
MvYnHb2uSnBA/JWGEklK/BMVuvuBBUAQNjeylvBAocIhlqlH4F7MI45ltut3v5L8
hVkWpk1lSslMaRD+9NS+AGhcixAHuX+CUzMVKAzVvnT/MB7gYPrv7YcuxibiWkP1
LCx/IDI6wFyzqRk2Oy86PFRKJxM3FTFkKtCl/zXeJNv+aYPqZ5mfNvk8UVVo92SH
sdkFtm0nyxYWRQ92GpzRGvOttBimsP+NsChhVZ6/uIEM13tjcJLZxun+lxXI4WYc
KCznAw5bzFJdwwNqEuKotgC9EzFFhLQ0fc5B6Maj6RHLqFpcIrveJ73bY76M4Oxs
vvLBNLAv6JPtANgu6hP+Tx/mL/9K32owyyIu4+PTJVyJTq/hXjo1V5olI1G/6qY+
C+3pd3G/sefv5zWRaFcotemKhhW2dQX4e89/JlGvburJHkogrE7gOZjFUY5c+QnB
wkMWcPs96CMh2/94Ife9sYCuLN2axWzKxv1bV/in9QofwSZnLKSgcdulY5mADURw
UoQObWkSwfRs0gBcg0BgT1qnXpovNIsi2ljQGCQRLWA/2LZg58mx43Zq1Mv6gyWc
s/keDDPBN35sF8RANfpGRIjCVK4QyWFSPfzxj1IVtTTw+dKKQ1xME8pDNkph7LlH
Aev45iMFiHCoDJyF/PEnsfm5r2h9fqnWYEU0MJuPZ2u+ZzOg/0N/qX/rqcEL0Jaj
yW3T1u+yMvylBdMAbdBh12azMYzHsWWs1UNtYV2/7IDtw1hl3SGYwXUUdPTz88+c
w2Oae78UqVGu8AbTFnyXBKwW9tXFrkxUek20rWlCUx1PiURXD/FaiV5WIuLaVJKq
cVsQ4LZj5SZsl5Nq+FFUPFN1uxUuAxS6MVlHwm8ytnfy+aw0yqr3XXYin6uYqyg9
DYEDthUVsPRUbmMAApfWiepjxilAPjEAzvrvL3U22TABwwHBTaq+LLjZX92LMsXH
A9CfzaRGoN7vtiOOnuiCbc2mCn2qXeJ6oyEPOuO1cTFuYQjHycpqn3AHG4/qHlXJ
pofvKQpEIVdU1RdXuydQ+5FHwc++B2RQ9QknJO4kZz6jva5Q7p5r60IGIRe+oam1
u/UTQXcNWK7pCXVMGngQ2fOYwqqF+32T/nlesSI14ZgQsgjusWGMUv1yd/3NiM1g
gmXzeZOzuymV8szX54lb9lhMXyT7ekXiNKM2RJalfrUxuaz2Adk5OvV1zuZriI+V
bcNhuIS9RK+tEY9E1Wdkfjddf1cOA0g+IL22MnuOJz1/l6WH3Lhx6qcwo2m+Z9hP
15q5b+LeZ5SHVSy8SLI/MaSRsQV30AkvAsxCxO7lFsyzqbM2umx31thQEQLziv5e
x7+6T08ryhX38h57tL1Jlf1NcjndjnzjHTXbbyfrxJDMDEGISXQpS1VUWA9hcqVg
UkqzusGlsQr5YVI13VJiJsy8zxxuJQa1apMlzYzJ7bnUos5W7syBZ1hVRHHWI9aB
47U6b1yICo9NJtt9f6F6d31C+q6xfrSyGn94pge4qS1VpKAiaLMtV3+19ciLa0Is
qN0e6NqE9IUJ46Eyy/kunkiWzg6tNckGxnbTC3uT8gqdwOwR96yYWq7Vinm/44sw
Yo48T1AakpAqSa4o3hdp335x4DYUsZOaJS3X3Oj+H4E/p/wBb1hbbZ/OktJnOuWv
GectQ503mp0zHepfGvmn1LWAe3Y98PVqr5O5i0ADXKAMgwWFRQRTOLNzW4RTB8UY
fAsT1ud0V6H8POoPqLMMVm+Okr20yld/UKO8bJbdfjAg6ESySwovr3kzrzAOifbj
I71eNifOx5I0x6AttQjUXmkhY1xhcIp031lgxNhpa/hEd+55CtFCd+XgjAGgJP6P
6QBOncBcFyjLIEHgKadLUa+FIgdRI3T++QEL4wv1qFV92Xhpx8gov4OKbrc7Rj1L
UgSjrp4rMD+wRvdTE2DX+r9RMfGJjf7t0AJZ4TQxU8BNam2zUzbQML2HzuUx5vGD
noL3uF4VA67UNGSog40MgNeXA43Juoyp2Ix3RQlDzgM7J4BfRjQ04lq5VMnXU4Bn
Y0+ndQ3e4VZwlVLE+M9rMyanGfkEvTUlbb3RUvpxoMy8IdNzxMqgO9j3QCmGwJnj
savpotVbEg4Ej0ZSpmV4SjQ1kq4y1dX6+/kj+vK4TLgf/KsA99PnlHJEBdNOJ5oO
ICkBAjH1jfNmqsXGUGxdLjH85h2jr3EGaYXQvH++R78kNiqogL+1GO7vY7SppOrx
GuoMuNXCpqiXWpxW49+AQ5HnLbzbXoXVyMhq+Erq6GHeSgwLPF9bIoDJ+MK/l7Ie
56H2fvFM7ynBE7xqbuCv9giJtBiYfx379OvegUNAf5H+o1OiyFWFlEigX1CiPyCO
T7KAAisf9V4dOYWQQo2TAx7oy6eMO+EnNIzk1H8np1T/nrGNB/j22CqP3SK+fuKX
HkQNaybyQXaormkFg4p/ktvUJt+MRAXEwN0fJXLhzswvYOmnEuALr/NA/OmZhj+d
x3ymW4rRFrcz5fe4QQsmR8EQQNRX0gDcmKNmgbugLv+FUBpJVhQlvJJtCj40qbyT
82IQu6Qwdq+4A/nM+ZNv752I8ZSw0kpakBCecCw4Wxo2PsIFO/bw7bRnCz/2FDQu
o6+kGpuV9qaTyNWE8JpOJ/0Zv/j/pZpT7ZJ0pFQAilTAYV1GeTHXrkv6ck1ay5wd
4TEBCLhqmfIZB9XgfPEC1KfuuT0oTOgzzRxcbV5mfV6rbZqcpJaFO7gJDTVkz4Qt
X0IM2HFvrExHNgpE0+YbZqcVdf/D+mps9sknGP/Lc0ROI5GB5U3nkN2DGAMr4knA
GIs1RBWEobjaNNmWazZcSCKHkk1wl43va175Ix6g9ndEeraKi6rQSTWqhhvmter+
xOgsc4fzX66DTDHr1a5wp1QGAosg2TZkZPCQqMetRXIeNX3A7Gcf4iR6w2E5gqia
MfLJr+iYXjvx/xg+wew3TEcxliYJ5VpEWvjPamAwO04X5NEJRPeCSgG1dOk9gCyj
KnLPgQAIj9uv0OFCmR3ytaGGNkCiwo+97h0ar011burhder2YB95v6UOwf1vKbNN
2jDyGw2ZKwcAMMlq8xXra323wEAI0+XSJ72nhDH9mPq5CXn+R+NHqF5vK4hbrm3/
Zi6rZOKeahjz2GwDXaN5OOfY++Rr+Ks6y+kRkxEzjLUr5MyYKwiJeuyWaotDyzQJ
4/9nRu0NyWePH9z60nNqKVilGv8fPuTOiF439f/HCFtu9+qOcp1Q1icZtI5dkc3d
rGP96kFUGuaH83R8F7Yxyed0s3+GAuEhaNfjQg5ZAhhJ5C6IOhqVP8fX1egXNEVp
jltj9OR3mRZFBD1aT0H1ClShEhWgYZseG3PcpM/GyVwuJ1jlVsK3PYs8SFKOeRxG
NP51qE916HHH5e/RnKQshX9t5mueaTOBHnqie7cj5zXjmWkZTNX1xegi1IK6+RWx
3gqqItwPKySpTrNJtskXNrhPatsV+WjnUZToNyZ289E48TA136PZ0n7YERTqvVvl
ZT2K82KduheHxP8zMDbfqBkQzujVdq/Z6hJC+3lUuthWwmqoiruLUaOhMmaKHPVV
EFm//7FmZzsv7gcVNcZwa/Z8JlmIxza5Abpbb/Of84TySeUNoJOHWC17y5uL8Skl
tnaQ7JfKzVpZo+DW7P4uyRgchyw2KVD5t2CdLzDjFu6itr9kzVKFZ1NdRpLsbuup
WOf1zwNp0t/KgHVuiI4Ubq52t45/xkJNy0IDs9ChtXvBe8ayCjI6SZE+kJGDWdy2
nVbuXJihseGObViIa7vGI61JVtufhIwzuGV/zM1vQYQfl6FBDGWDB4VExrLNJKNa
OOxEYwqoIohdx85d0ivAxp1N8UYlv9yjVp0WyEWe2NfBONwiTs1CsbJ2sV5/4FTD
cwtt86fvfKgxPLOqUzNmqXJlyWjQVulf/M1Q48xUVE4RdQpJ6Mfk9D3vN5Q+PyDp
yG+tE2+CSLLKv19MAZpgzYA8KH+tE9Z/dFHPOi2lJOnyLS8tuafsbiPLspL3j4v7
kGCRNZYJi3TdOuinxvi6spUpE787gaaap/vkYVtzYjheZNj+yYXNvZ1BXZbHQp/r
OiNy/9J1o5xpLZP/eGzL9ucPQTcYIoxm5/ndvSLwH71qPF4znYAS5UV7ts8uqU3q
7nQPRpFOtk+mRVJN5M16agN049sDd70gxsJJgTNneMB0AcTclgDgOgjkDLu3pkD9
xrTKOs44J7RTGRHtxDfJNF0Eeheb2ctzCLDCI2JE0EM4iU1em2AtDPPFYhDzOcfe
xZE9LvKrXLZ3C6OE+OmBT/GuRetoypyV6amIFYB1xYgX/OOO4t9Fvyfi0IIXxRph
xnKuHRQpOP/qXJhYtjnXsxXfl06TlNJ9CkTvdKzY/LcnYmZ55NiopMgN1bcpalco
DkCZ87kllctiYembrdA4kuLV03smcKDQmJLmfMuQbtary0NfMtjqBimM60WAIFgs
WDlEQsJCyywl6M1iDoQK3tG+kat06UCWD5CtZiC7H7I7cXyFpms3Tq5wv+Ic+Q/k
Cc9TtTb1F9RIgFzfT8bhY8kUlmZtSjEVfJKJbCTUutsD17Ny7TWgfF5P3HbD+gst
o7tEoBfsIJoRVen2JIX0oFZpN3N7oh/C2V1c5U+Z2bJjAwNklqewSAx0VdBe3yE8
Xv8ytwFA29mb4yGdrTCprBGV/WbcWiZNfUGzSyTJurYWGvJoiYET4VN3mMD6NojT
wGwM8fPAgudYP+5TUDnJskwv+BMmHoR7pAcPNBXUZ5GuOYRYwgTAXiiJ67hFxNnh
h33M/js0XJdKx+eX+cJ1wmvZkELKgKkc2tziPIxl8HDNopglSBMZhjY/Gfr0JISF
iyR1JHMTonsN+Sc4cUhYs65+gm8g7MqwEEyuy7N5FUbX3QyBUZNGEamO2LKTsJXF
gXhceiyrfgTgXLZBct4G1C1lRPO01CWtTUCjpqY6YBZQa+o/aKVdXy4WpqIorWyt
Mg1NaemVEsngZE7XYzg6iEV6IXTXbCJgBCdRSYsOnkHpJ2R/eoN3GzBsf2W6sj0E
Hgg/O2zeNLOiEtKSuxd6ORsrTULyHowuyabunBN9N4PhTC+DS+BjqMgnQW3iVvVx
H5iiRwxjLke5XRYCw/xvtdLmI90UT82N/O4fbSb2bASUHdwnYQzqUSvYNqUwCdHh
nrmOffZFCOIYLgfK4cX0XqgjSq6XK+oiPws1MnXuHjkJEihBsVFvLZCZFPeQAatX
jnnvnbZvjQzXl2TCseBqEcK0WISI/Vv6irHuD2ZJT80NmDAprO0QR+JH9irYungG
+8ufu/XL8QNO7XMiqN0tE0Aj/A7rrJmtiWW1r1VlrglcJnNr9GrgSLGMkvZeC2MB
rxY30y5M+4Pw8Yuqs9DxqQQVXS5TGKMeQACRRB0CGniVqmIDTwsLmwbBcOMTtiX1
YXV6iEqFDZRTbHBziOB8RCS4UGg8RqeTCT8iYwQURMXro+EybMVPUA80PQiJ3Uwu
ccrjMLNveGQ+1aLkM0mDEmbmq83i3BmOh2yPG09HGvLZSquO3ktFU9aP5tE0gyaN
aWTWkEW71eJsXZwrX/clLuMBPL5Km3V80/uY4j7wqwFVvWxa2hmway8UOQKQGdqn
13odhCKf4qkrPQck+c1H2UDmKMIR7TWZ4qJM5jMkIvtWhY3O0Uzv9rE//YI3oZp4
EyNKhysa0tQMrWZHNhAnT239nuV1ExHfbSKNss+F0AcStIdc6m45kGlQqKRZQTjF
30lII/4ffspwQNiBQ2zJP0DUw9mC3SLPvGI3uJC08PHvWjn1bISu94i025gmqQ+9
/LSpHm+hxxQ/gNtKYF0cFEvZPZuTWYQgYw3K3VVDH0K4/U0kpowsKlgH5q1+pMXG
SIWWiECIoaNLmeimKS0NbC6DnPv/mblxffQPTHw/wAc54rxzTFoAXa1nfg4WI+w1
I1tFwVVfAtRDNHIhHcdQ4kB9cV0I7vnuPGgemFmXXEJZJDg0yKlB5YxrIjVzO1vM
djbkQJoFcXLdwgNTksP9IJOy9jhHWchkSX5PmbY6XlNqq1Op5P+K1x0Gs9W61qzj
0yfQyiCPcbd/aw0PxDb7MD7U1PYafdIIUgD6Do0IBYCwvmEat57bgONIkRrNBwUL
1gLftHR/sVpi6bVkxM162MeKzzo6ql4WiXs5g/ct9mlFnOAfNa9yRXR5GAupK3HZ
iQnbHX7UVqzqXEhC627+9x1WxxWrOfOfzcovaeGS/nz0SXnapGdpnyGAU73UKqy9
ojwZSISjyn2kkOlY6t6lk/FBtAXl8i03M8sQcUgN0hxOkOLwbSJBnzC7S8rb1KFZ
wAA5MhVGo1PyjEF1D2xflO18yAsbrkoEqzXCHMojreHHgufzuHstOq4DwGHfxSju
o82mxPzR5vDC1HdU1lVvAOX7Dit7CgfpI9CYk7qK7/wt/kRkvKLjfhoFjRWy18Su
lHzSOkKT8NIHdTOrA4+/ryPRhIz4a+tYMAaD6Ljo81IHnIh0fhSa/9F9EEFV8o6z
wWaT7BXOfGnubEmntcgHSMTLRWrK2ssknQTx1UybqPEmFwHPhp6BpvFRgT/0h0wf
KEuy/IgZo0Oo4zOXpUxNAI5yXlL57eMMBCOBwepyPJ1UDcaxjyzDTnlqnqL40f6X
1ayhczZQGzZnR9g1x5HoE8BWC8D3jlA7rXa7uVpQXfQq7VWqfT3ya297nLznW7At
zVUkoAOmPNJqxigDoj4BR8kNr3zMbf27nPtTm11jXVd3B/NkYFgk1upCmP69nlVX
Z93olRT76jSJSfMGUpQbpip07TEWKIl4fp9VjPfRdZA5Gw/UtHdBOyP/CueeSlCY
7VuYXBUzgOJG8ssr/GITVbypq/duyCiFTL/HclBlqainPT8r7wRG5+4Gu3MEohuh
GAbfoo4etwLKCxyRkvHI/G4wudQr7/A7OHsZIfuIa0UXESV3WSp7FORdkQzJydRr
ioF2ejy3HHofnxWtDOp5Ht249LsIVapDL2W/e3DaOo0mP5pYPRIvBiFGeW6APcNb
0OrAAsNGeKGFFJpsTN0zkpPahhACsWE/MB6zZgC5JLZ7uvw6yc2KaWtSHxYIM9HP
EoH6PvuJ9/bOCZiw/q4gw/KJjEx6qrPmIAg8Wyjw6mxYzqJjCtsvdu75/GZJOl/O
qsCFohejsrCVaQO0l63OYFN3QuwfqajWNUYVcFl+ZahKTQL29HdE+7DYbwOHpRdP
EdFs7waim0PsvBmjxtr8KVG1jYwgtgprz25TRPw80cNXhs6s21wknLU0iC0o0J75
dLcDO/iVuYIxoHNf6Qiy5JwthtEjx2bWKQ4O770K2i/rM+S3sMfHNw6ZA6Q6Rqz3
AJwy69K0Av1y51pv3PXgIlp9mazfS2ibDCcVoIOTaE/cOSF4UDkL3f/WG3xIVKRL
tQfpgQ3p7bo0mmnkNLRLHuoZ12LErhO19240mvdUEl8dLiSytWiai6gmCYZ+EfiI
5AfC9TiBB3pKPd+HG9WVbHQatgJoalrZSzfFd9tx+sTMLfl3DNvpW2P3C/VZ1xR0
hNs3esUmovfLJjr4odIcxWDLQdQI/dZxto0LbD/tsTtNOybvduaI/XCi67BwO4tq
0u6oHUlThRLwnrdG0KKYMdV90Q0Hyo4XCPXH+biFCANxdgD8wd7yiHOZeXp5kklA
zhI2poqCKOqbYUGZzrRozuGGwaZoihwSxtYT7EKrTNoF1dPihpg0CT7AjKwdxk0B
127AOqKjHYsjyr0m/ahyZHp39Uyk7jRkIhWY/rJ7D8akMKkmYB6xDQOiLlcaMXhG
xOmt2C3KMdiYMzBx3To2QSl2yck0m4/WGPhgln2yZz1ja46JXM1xAZdWsZiGAqgH
M7rkMd7pkyZXUimcICHofWfL9wv7d5mrL9XeoWvW2ImjhC82fVT6hJj0+lbc5ICt
w7A0nl71TEptXb3nFgupVfmXhCbaBG/2omjFDA1QdP4HDClQSBe4fc8eaw9w2OM4
4pC1wBkrS3Vf8vOSwQSdhGgAJ9heIx+Nw6OmWtEKOrhBvZQ5fv006h4/Aig4v6Fd
f/RCG1pb06m+7WT6yG+jAjxogUuTNCHDXiLWJX0AbXjFvb4eCloQnA2GsL4rKDdB
skafnGtrd1RISZ7sFhvQ4WsydB2orjAJcMyoiU9RCFOlnN4FM5usCAJssuL5NT6s
VwFrX9krLshQpwXrVBiAqXRcM0kVA8F0iUGn8l9kiEfuPgmOqCJ38i+OigBHlata
nJ94AfG+ydOYyRkjW8AxfzNvJl1rz3X02/ui7YgocZw9fD4Hqdh88njbtGAt/ylu
kRMvaQ0/1TtfVRko3GevTetJJCCUiSIx5AaQcr3qucliXnGAXZTUn9fc7HD7IjlN
vwSIAk8UIK3A8p290bNy1gD8SLvmlxxxJFQD0rL7MrYen5LIFOBCWHr4toxlIGUl
8yQhrJewO7GAcbDY5NZmO0AMHuWHo0pH12q1NNA1TkbwZO/5oOyniY72RVvHRg3+
5+PBaFZOZwt7i/6myddHfJDO+UtKBWN/OGcbxHTtiEnozXJlvf/QmvCdVvKooyXy
p/Oq8AXMpBhgbmZlZ97ZdW0ZTTvV91wPa4NvbdynHX3v8bghhRRupJ5pDtuWNCEx
oVhZyY8ESivQ5G80aJjjxoxD41uoUz3JOqQiDz96VIiHLtY1EkwWN6laQI5zfcbI
2MrbHOskiom/DnACgLs7IT1GNU+AnM9lBg3mhWn+1AA4Nf0Y4SH6SAStfl8hp0k7
ST4XoiYe20jw9L5Ym25pQB4xSplrXBif4dCbox9IK1N0NKehPLLXWlOqk6JuA/G4
RZVpyFFuLtB4qRUdX9KPgEVIyy0trwY3ZamL3yrZKJlVQgyQWD0IQ1LEPrOnKtCN
eZ1iM+THBhXe/+SLuIroVD1eobuv4vje1w7p7QjSxo2k57MolIlEMt0pfu0D5ppZ
XvIvo+xUxQtxgZFzNu5+licvNal4JrTi74OKp3Ja2gsh6r+kLYgpgesYt3dksS76
jPEGKqzhmDy6sD4tIcmwC9W2uNbkHCv44BFm+P8S2DcBuWxADVW3fEIgzxOOZb5F
2aY1akUklcKRKyC91RSAXgIWrjAUjHrDxIPuHoiKI2Ar63cXfDgPsdRk8xqMJ5X1
uRHy97346oKArAzUEStg+lZLH+rlE87/pfTUZDkTDq/a2uYKe5iZGQWFEeEfBWMB
gWKOE+0hKGmSUCKMu3zPjR5G1Mq6dvFrl/TDxdCDIFIyouv7Zq04MXjHCxr4gsFE
CyeD0zd3jVk5a96DFRnbk56AJFBEdSAP4e/SP/jXGXt80JiGlYuzrcUQOiBIjIy8
jTOhsrOinD2YWekgY5NL6faTlyEei4eonSwo8AhIxY8z3+ZluQwKBD7+Cb7Iv7x/
9T5QTdPyIYjPf29rPurcDx8m8JYBS9dKvwNdJFupbgIAG6CTLqrCxigjihEWl9Le
dlhe8tufSzGDVk9l0QQAjbxQJTUmsXHX320lZBKE1hvWgZnQQPb9BZGMMIeKuDR8
PH9SpH/lR2iTPmbB+fQETmv6cBFSliI5734DXjMpUCeiWpTfemyDNyt+jiQuhR4x
i9BafYfJChaqoj6rJ7XXLHn9Blyy2FloAGoYZ44ghsTixyJeq0TSGl5Ij149tQb4
U9EEXqSNAv8hiRPmS5ncXSZyuIXravXWmUVIefRo+JfgcvrWKfCtxnL80Fx3ccCP
WF02okT3hThjXaXZEsYsWrj6tcQuLkYZFjiHtOQBA9ojTJ/C2Gat364WdOzw+DFh
VktQxng9Yh9HPBesNFba5tQR3XjRO8QtGzuDJ1IZ9euhT9mUnMSSJOgKSLWN+aqU
FbXu+ndcN12YmlnUnOYYg6pq9lC8GnykjPF0WDGPRCBtx/JVRe8KySfqErK9xJUN
kg1Rzcq1u6bK+Qgu9gXNqVUGChxLUPgcGTvSjgw25pK9TAdu/F7wTIkruBsKkMsa
S0jGeuopgkcGXlU0DvOiUCN1JDqi3k55+m3MAGpN9gbslFEgqsvDPTe97bCz8UW3
q68eBxKRS0NI7lJ7u7W/weCa4mNv10qRPZLiG7VnBu7dZ/WA83jSJLJnR+91Cq34
BvqPq6dgKDDNimxKaEMITwuZuBolO9Q1TBuyvU6OI87gSUGK6WOLA4QVzJNKx2aG
TE4+NkR7I5HKkdoA3VHzVSbKKtlysbX0PwAxA7GQpe1+BfSZmeYFDnjRLo+kY4my
+dSD5g1/QqBTmgFu63+FJpMugUPq1gXdeSm06Wm5wvvO3E9Oz4F7M/NEfnt9tzS8
NddNWHmoz/ApQIxmuR+HJ4sb0ZTX4jntaFERNRLWMCgxAndjz0OiNdHVRmd6w6dv
r0S52jTAKU09NFJYdE5t/CEyChGaMs9OU19ftJQD+MDW/anSQV9qR/aVfEvGCzrP
/K+Opvp1H1ud3ft7P7J8zvrIXxgezvi+SA9YDvX3whGhvYMpv0lpGTXDUiXiTy0b
OGXa+9YEkp8s+mcxVW7Q+RvVX9CLh+/JOgiRBG8bRj9iUPh8uPiE/eQnbvHCRQjq
QrALkK1scWr5m1FBq3Go72t23IBzFKg9/8JO6VZHZAUpoIcZ54MohzCjSNlUm3xs
+Ms9ujn5OPzU79KmVb80dQhOcvWi3CipUwmUroUym/pQ/Po52NxfggJGtviB3lXg
8c0xuQ5gzZma5NGG5V6YpAv5nbk/zjiWMl01Jsa2foNI8KT0GpZZulHKZGjSeTtP
Nh8bFTbQgp011EbZZwP+VNNDT2K1rF8NGzvcq/vpEkm3CS/IBqj8dxhEjIpPSftK
OCnjkvjZVSpgEoOwQBEg8sW31zy8T+SSidzYvzs5DsyQxD5jfenST7IiheQfLzo0
KEs1oMbrLB+jpAVUb7xtW89besOrFqQclUl+QC5axMth9mfxukWmA0g+TAtsGxzi
8KT7vXUQaryp5dukr4HjVKREkWhuyQ1ME8qnAwWptezKZQDMbScdFLskA/fjoYSS
sBGkvALRzQD9c1KJkU0pQjePKwBGyRSIdkFR1z01IiTBE/GDyh1SI1Io25HMzXey
jJEHnQu10KEr4N/Jus2U0MB8heAeWWTYEolcK3FVPDFkZ5T5+NGPK0GFb1Gi4xp9
IGfn8mbOW+uu+F0jQT/cDbVAtbXV7bO0JMB8zbem/LksYes7lHgS+FTdjJi5CKD3
vn9rKMsxHqeFJ4G4kU3VkvEU/7ekYCdOxs32w1uP0D8lp46Iko6wZgb8QZts1yDm
K6SXxMQ3dLOLtm621pwocsOT/GuXQ283j/vYPtnqWPwXc3jZjVogozsgfbfida18
tZ73Agw2hyNu1PfRIa3Rdbi5Cfm8i5p43WvasVbeLaJw6YU6eTILAJDXg25NhpAo
emNVydjRtYTjRUqu+TkXeXDP50SZv6NR8HRYh/XsASu9JBPzaAxbb5uS8mX24+qE
mGbTBtQty8vrAHeALpkDDjXzUyKu4ZmdA61Y0RDgZLpBvXwxNH+s/TeC+MPvK7G/
rNTPj2ac7wQ/vziY0bWGfCp/dwI9BVWh2eDQuRUfTCmivW1u/RLbL0VpjQEKyoG0
XTsoRwTTwdSvA2dYd9qZ9O9f9nR75LIMOlv37+BeEZHt2pX+CFx4VmdG7qFZbjcl
NRNdzTaPUkn+A9xYIaFCkdnYg5MikTJeP30zglzOO+H0L9udjDxEWv/FEF1GOZdb
igryciwxSbVKJ1nrmmOckbihe/Y6YGqkDxoFrxUiG7VmIu2zbb02kNJLS8t4z8Z8
WMI2thnHlmFmG6GbToDt5u7U1Uw41jHu/ZkIZYhKLUZ76IKD0MTfWhNWGYOZmtg2
Mg/AXFe++vtpszj0f+v2+2wTgUWdTnJcIrCsKS7kxc42MUegF6bTdfD8eaVM1Whs
0j3S3Hw87B0i8NJDkuG6p5TI3gcXUrwoe1DkRhIMJQmAYsfTh1S94FYFjpBp9h29
QjiKiy8em6g5YKqu2ET6S5bD4GoE9UObX41pe7s/kHnKS0jajyt8BDLBDfdFrGKE
4QozrQWB3vLptzQIP8/8tUOykwLpX7geBabZUAKFwpGidsakSd8gr5IivICbK4u4
tvNe7hmdN4x5N0YNyKzM8QIki1/Yq+Qv8LZXnqlX+1LXpY4ua+ANaKUkOQDI7bbC
GNvXvII7YhvHyyEcvvk2ORBreWQut5pgb7+I+8rI6htN8IAOKdihdMHozn/6DKY9
LbsZTWjWEBqbIxz4FJpSAMflqxiN9nfmJA3V71HX01a91yms6wlPDlpZUpnqclZC
WU5+CADxE9GmnqlbvPeRFssN44EodzYZbntQmFAZJrlgsWPbX7MHgLTg3L3oW3Q+
n+QcYdRontMzs/2i97jLi92WBe82Ri5kSgeEZiOG6txsWIJ8s3u3PO2LSFJiYj9z
fdTFv+DageV86TM4l68nrKTy77fZY7QBQptRILUAfdefRW4E+2lBgjuLT11WP4xD
0HvsFLEIArKO+tQMxkryZKqlU1MFGys9YTI6Uvj7+IuYQvf5kd2hAYQMxsw56Nwl
frTa1L7SBjdzbtTU0da/qUDWs8e7Zq3KS5CMkFtfky5N230FFKkThbWbdDD2LnW8
GLu7Sycjl++EM7ZnfkhPO1sjPS72qXXoaBcu1bkeinF9qWQChf2ZViNAN+5gClB4
vnJMMPGF5pX1KCgpB2a30zlpdGHFCDxWZVSvAOEmurGsN9FGpIM474NDg+l3kg8m
hAifHWFmjaEyZFq5kJWDcXQ9pPe3ynlE6lxqR33QwsmbME9xJWrNDuOKeWuPLnQ4
NwVWrfna6EqxIzmxzKhAAPsmE8QQpxyLWsFjtULoL+iYqIa681TIMRAqExkxwlJz
egrX2lMJgtSUFSzKhFOL8qM+IRp8eIISZnO+PiyUcYAwdZqj3pulxG44s1f2Jg+7
NbzIP9o0O8FxabLFrQt+/vaS5Wx8NhzA/0pyar7oXFLRdQqWhOCM2t3r6c+RU9f0
KicX41xbwqt0/6+cYKZcGowxoJP0b2GSljqB+onOsi0b4HE1cQ6qhwQwVXO9pu3k
JSV1W/mysd1GmoaSyEMem2aKhXPia54QIFg0hcjz4t/YqaOOKKjTK1dtvYDh1vki
Chwwq4gm6xqJdH1Scu4KAjlse/UgSWdHvC7Es+JG/T0ayLvbGrmjmLTtAf1Gv3kN
qbQldkYwG8lZB7LUme59w6YVQjH1WMwW1cEWzDjNlPNi0fVp6s4Ar0PsOvb++LP/
J7GsbAvYkSYmISKQFGvb+CEUdcH4G8TOwzhUkei4SmZSQLD2qHQPZ3IBgqzYPwBr
Y2N4b0aQ2ZAWs8+52Ks3YgyvNtexa8bFASAuqYh6xx76BBYvuSRTYH+cGZumGHiX
Jz5H8t5P97TTCo2pojROBVymjCjSBBH/GoIpWZovY9wziISTl7Z0ueuKy3Zp5mhV
Ou0gkeymWVv5vZeVFLJ3GgdjlUvR6lHQUiul7CVk3NTWJbannyDdCVAXg5+ytBap
lCQW3W0Wol/AgYNMygFST67BgS7vD6Vke4p2Nq34gFnE6tXp8oTSAl9wBMoXahJy
L2rtS+U/7XMtMLtLLHlBouMZOTBdjqQy/wdN+e3JlSMEUyl4E8m4zSoIYISq1fQw
WSbOu/Wz/vsofDVZvNb6tk+wvCPkDvnYAYLI2zXcw4v1njTaBmiQCTDj5tOlBaLg
eXzE27Z41LwtD0wKfban4UiFi5s682yciPNk1TTxgThheKx28B863isCduInDEnU
I438fuRX5WueZVMTt4GUpbL92druWU8kfJFj6bsvdkiCBlYjdEiPnYAiO0tvV5S1
4t//YibmlQhhO9Y+Wo158y3KvrnZzzFy6MSiqPYBBYmLKFltOFwfMRtVDTNIG78S
PwpG2El5abkHawoAdiScpQspjMJznTdVvN8rWT2mr1/vjKQs5jBoV3l9JsdZMpbs
REa2Qg/xinF09rXLSQ9sNZFz+HV+4ESUD8jCc3mQ1HqE9p4fP5Pzk13n6X+iPOFV
AEFavSH9H2U5UYs5/pjtWYxGJyXixe+a7Prx2QtTT64oG+X6Xa4qcYK9u3uOaaqb
aU3X0xN7pSTRTUxc17hVJB3FEBvf/yNFzG6FBp1u2ijkB5B68hbA/BTFctZ9eq63
T1muvJWnW+idFqa9U0uuNw28tFbjqKEtk2BHTWM8vprBD85velkjQyMdZh4nncCb
L0HQ52q6Hxd/pEClSdsxLqYfFOY9kzRuvRyK+T04p9oYI6UOtADVAn02EXz1QcYv
FH1+BUF0gFeo//Ym04wCusJV2YhEz7bEnN9Ty35EOItJMuost022aD7//U4Au1Df
fjv99kzTTRb2IfsgrWp69qisVdVJCLpQ+TkRDAbtjBkaumAHY2s05Hj9Od2R7oGH
GF/nfhhT6N8HfJo71Ws+uTW4ykVnyTeiMm2Orq9y4vDgXCDuMGAKxigq5KJX0g0d
jhk1U+wLmxEXtjDPlLrpao6DQarAR8nJvAPjjCnLr5NOxqrZhgOBzaG8oVLb6EOF
PLbvNE4W8TWfFOJehBngT6SlDA0mEWGe6fsZmu0vrKjbSH3CRivbvNYuNbix/IHQ
RIH5l/07nA3T3+4eW+/0zRXGGAbpjXq5ITRfTTCAgtFDWl+YjRvvM8skR+R4aBla
/cfoSpm5IDtpBrf3HLAnu/PP3RJoNMMQnS6bwXOWquAQRIfTcsPP1poqtTvRi6ZO
aCUmsCiTjGVNuHvGEijHdYvC/gB8ZQqv+4nNUGdtSDPsouZR+KZnoL1pB3ItNdzC
V56sMje+L58chqrNnHRGpDPI7njaupZ0qmOugORTWZn3+XiwgyHFMlRJZSufqicR
96roT6T3ZbD/2qLQxDiDRUtwL2uVT7vTsUnfTR6MAqBrpQ+oNxlX3+v5bVLc3339
7ljmAJBV9wuAGpFgmWv1mIw/1LaMR5yBKyK0D+OpPxaiuwz8QqRbtq8/t4hxBelw
tiX3iuisFONMP9gSn43KJsSai0zVi5+g1Z9KvIhGts9QlsV2d/UPGU9rOVkEjVIH
r7vkVXzSUElWT8tsDOJ4C4KAkxljOH5kyx94iwY5Gd3MnjOSO+qHJlHKxVkhGezk
V8YhuQ2TJXAv2OOdcKTVJS70aQfYxvMBj7jO84YEYZfH/yiGjl6Q0OQjeZSvfYEi
nl1kQGO5ltkhxixeFCoXbffadWt3GN7d1Nv0oypMzOrgn+RVCnLBk3uvc9jvBwG3
Mvr0Fs7yN3gEwMZoL1glvORd22cvP9OTFxdGbFkbEo7XxNK1IgJPQlSmdZVZ/yV9
5Zx7VYuRTlY67wlzsMnHSCuTjnJbds+c91ieHsB83hAkrpGfdrhDcwPxcvlwmfO+
tWHvXrSWaW9oXj74a0PPcKwGOteBb8/Iy0H53R3mmv3RfRaStjQGSuJYfkakfLg/
9WdLN2bRoW53DiZavEiPkkLCcgpKhOzeVayca6Dui69HNr3nn2amkiTzoTMckaC+
irQy3+4cNV74KuMbxhqhoTtPKrAkEQwEnDnftB3G7tI6GPUchoBbM5ggdmSliD6O
8jGzZU8IYRpTnN9yuu5aF+FwXKHcTEWhzFyO7WY0q5X99MbDZpiEBMGn114UN422
J1AWGY2Y3+WzExmJpHMB83yDXdZTZU7yToh8Zo33qISqKeSYhDTrSNVpgq8LiVpv
kl0e2OgOtCDTSAFoeMAgETx+I+CANe6Pu7yzS0oNlOqw1oLzjCzizf4BjErSwa7G
dU1a+W/4riNCOcltryTWTT2u3lGCBYDx/3Pcrd6d5J6v94VBjaWvAt9zwkWtOq8+
74beCr5AdkyXE375uwFC4usF3Gy9qGbB9hTEIDvGKs7gV30rltaeIRAZYL9tPb6B
dksENkOxXybBWWy9hS130jhg3WW0K+PzEJMiuWW6Xnm344PopnK3vHOcN67rwpj7
rrHhXMushZqES2J31kiHLQAKE41iIKbmhPKqJJLZIgX5OwFKuPbiSfat4ZQk1E3o
HCa8yZxMlI65jm6gcJHlcHwnKUVIaGr99zwQB2FaCpNVsQRV3m+GbxS0VhYwV4Q8
Rw+cFipzlwmH+E5nVYzV4nZMIJhDbn/Q74T0T+1mCJcyujPSnxB+iDPs6zoKdvst
A9/GpMgUKPDzmuz9kr5CDEFp3huQdo63C0EDWj6SdQveL3Hw0BKTbJxw9P5Ytj8f
+X5mJJ31rwsGbVgnDYBiF57tYpzUF4wS02TGiobAGGlX6nrVY/q1AYH8u0+FCYkW
5yXznL5Px6+65JYLoa9OgNYGoNjgowj71odORTTZ3vK6Y87w2PJe6JMD04Cx01jd
H+4v65nFc8MCy/9YRW9i/Rh7qP+HhMC16/Sx9AzsgKYHkrltvBpwq2UFGiEdLr8m
VgV0UFAhkX/fKh/cL+SEJtqJXj6S94kiSU2Ql0FEjCmQ4pAnudHqNfxEs9oyTui4
txRPanZegOySyW5NxG2i/7GxO4L68r/FAUlPTEq1CW+v3pxc+t+Qgsmu3GWDCg0S
yRdAObGUpbTJuhrxt2KRE+N6+RbRteydmfxlbL59gX924A+Knz2CN6t/kwGQFBxX
wcpV85U2p4GQDqBkbIT+16rrXlAwYWJ9wd5iAtbrUvjBCrQOylaGETxWVK4/gllw
biROKodUSakXOlyyv/gLLyrfx5Uv8WirPe/ut7l0224gDTN51ow3iQ2gUnXRqZLt
p1EEHsASQ8IfZHOoMz8xJn9GT8cTG3owMD0kIQoJ61xPvWk79Rk6/hlHNZpl041l
qFlsNnyuWsMUOmQFA63GgLbnZG1WBn9VFcfqLYeVrEUb98NFjjCbUDpmoHQojPOb
+BwMrxCtgvPai42G439DjcKObHihlMi2834DWqO0PD4y18oW0zRZsito4B0X/NTN
aUwaz9GwbJ7Vr+0wSL7rjGoQAqh0x/sPoakdKyJsso/hi+/zkQL8tKroC0k6dixR
7MzeWSFwsLQaAZ2q5HxaClRfuHr8rKqFroqo1IKqgSzyhz56RzqeLnYGvLPE8Pne
xLLKANSkvy9vvOgq6n/WMvq15lUvkCb+XOUz2hyvtId4wHYKl/20dIOzACQGFzp+
o4VQs1UOwUmhr3HTFlA/qC7bJDWHsr0bfdi8BlUh45v6mWXjjNtQyUnBY9yH1/ky
o5WUgV70SlyLxrzD1PW8cGLaOUJRPsQZ4YIDg+VICHa4XMrsl6L6oeI7Ifc4GRJv
f0+lJQ2DMS1ccUwAAZ12x2KgTY7sFghNgWWKqcJfmBxm8FIEKJUhXe/XymXTxaCZ
41esDftd8RNnNSBH0zOBNO2iLEr/iU9WPQomZ96DRN4tlk1SzEElEf7l/Y/3ccgY
oQAhWwNAE5DloSGPNnEMKwOTS9Y8CejzyMMsZKg68hluPLcwfM3bSkL22LWOhMiS
fsCL4BxETgX0SCOtpdG3HOYAdoB7gwOPTXQ1g1W9LCe5gfxb6DNUfzNdb9Z9yPWH
wN/pgcQDvOCeC0ssQvhfIlhWqjtf/V8YAwTDMRj6NaWj30/TSkp5SO1F4JWjGCQ2
53CT8RShymVF+UQsGvvkI1X3aIh76VnSqnOHahI4QkfCkWHydvJEqvmAFkOCWSLt
0aoG+spAacK6m25KwyUTmLzFTcPvxnxKPjfOZw/Pc2JdJfoySeKfRx/xYjdK0XOF
K78j30+iIvNNWPCE9UvyZYfVYXHm5+osuLVBKiQHn3BK40ZGXtdyAzRVIGIYMS1s
lnhAlLP8a4W3iyO9GLlVdeNLLw9cvlcV7hX3K9RKlI3lYRoOCbWbD0KqNbwDhDwt
LO6YNGHXrm7Td/PwdegBkU1appybMAlrz8l91pIriuDBfefl9ZUVunvOlL0GWarN
Vmj/f3baarCbHejVFp3hCfXuFvzJqVeOPTIOEfXkAxNEbzuMdiZQ0QNmJSORXcvX
T07Yg7rB5mtAcVDbkXxUVbLK/xu6m4f7mb2FEkZmykn04TJrBwCq8qUoti92jsuk
VJB01PWncMj//BxKwvB96VhFy4EvSo2/G1wFry5BkSMmqEIO6AtPbjJLoDGDRfmX
QW9duFD8VONSXsVI4q+XHogcd4RktuL0hOfQs8WTwSgzLdpnstBor197HLo70zuo
9wsuHbgnDQi+uCYlK3+rJeTJLmg4J/ksCT5FOMQhEgPKkHt2L+l2sYwP0xMOZs/a
TA5LCz5sY8+5oXA6X2/B5oxqzEpzmNl+/xN3zEFnGqXXpYqNIrXOQRNxQ3V8FHGF
kAB/c0ww2Fstkrk2cVMRNXupEQZ7c7/smQyTUrzxNkMSu4LD/hen+J/+ZtkEgQJr
pJ43Dcm9WivvwfuvWzJZqlg6DIYulkZHp8nVsjdPuQVcafuOPPk5Ta6UPN7Jg0b4
QEtNqkvanPODGEYELRuyKq9TAlAuXMfXg7krVICHDw2Oqiq2l0KL4E/kpJp9cjLB
VWorSMzpOIIHQ6XQ/YuGk/gCPDPfhrCwWxwZKUG7hKB0KXRHNZrVgAYTX5+nYHdO
JKQaW0jvQ/7KdfUy2Mbid4OAqonUxagdHQUZ0OeDywf+5xhMHfgQ52o7EogZBHrv
pyjj7VUCtOOctAC305EmmfD8+zfRGZs6wuIVvUcwJDkB2E2K9ZChg9uZS41a7dLf
6TxtRv7/47VNtrnwJl4eLbJOtw5Fm+GFLglMrAJmzi1zRvaZuj9KPBHb8qm0aLf6
nZFgKdvGhGuI3h1Wx4hNlzCemet75pSryuK62mlbfhgnjmnyEzAtM/EqMRVz/S/o
mXfXJKcva2ui1SOh788Epl4+LHTuJ+/LRROMBdIpaj0z0zCZMPnMzrIlaj/WoOpO
syJHrS8f/jXgyiFDYH8tk50g7PrdFe51MY10nDE/h22pr9zZwPOypOKu/7Jxdm+b
d0dWuhupA78rXNP1lVNRZ8K+PE5DBlcQ0ZcVLG8Slwsb0PQt2fPWi3it9Y6tjSWm
VhwGTop4QSrkZlspzIW3vEvN53gYpiSvY1gpp9HsViuBeLkCJ4Q6UzOd/bfKfQ31
JggJhEHwpoCOyful43Ffh66o2saMDLc9zfB0v3LWQ8XX8uo9zdUa9GNeLl5uLqOX
Ca5GYdpFeuKML0FKaBBNAaTylrsxJ2AedfIpUC5zMobGgQGZNjB7oNV5wPAO/d+N
PZkku0gkI2PQ0tuNfvmV/lFgTfrBcCg6XOmaia0AtIQcKaVktX1Gp1I1Qui2NtHk
T4L0ptI9vw4+OcEEkWnfDxa8lhE1dRthTsYMX2er+w0NuGVSBvSlR1kWJNucF6a6
AExwWDjZogk23n7JvOaSKXwh/lARcBz2wyfGm+c+kYK4+Kp05EYH0R/vbPk2X/d9
qUpshX/aY4MwWZL2mS807i5ZIT1atwJKiqzyIIh4LR+9GUgqPQUJ6wzhuXZy97up
mRxyDTg6+OhwH02bAYvNHD0jBwELsEybGSyXfMW3z6/pHYJsJ5LTBUkiwaT65bcS
bwY1gi+8LeeVrT5c0H6b6u9GctxJLdTo7G1uUTI1kRB5RmVo/uaPVxoeVtZRxU1F
JUK9/FfHDlKQHCSIjkeIc1/aWs8QVEnZ3uIkqdvq76+cRMXAoHFBt/Qi5YPEhOca
oZkLH7B0gDMwQi26vYVIzo5YNdzHNTcIBnlo4Tag7AEHXmTZgUc0foD4iLzpXqel
w5wHMhdOaRph4fa5Vv4bJ8So7keYdVH/l9VIkZKF2YWOnocUNGYDLLcPOoFjUo51
qseBhAuTuzthMFvXm4fjWatRPHpiZmiFxxL7OMHPmYvmDIek58gSJjbk01Kor1MC
M2ENxfhw3gxpe0uaOXMpE+yOJskR3aq0yeVUtg2EiYpQYzFc/sV5y/gW2HOobLV9
dhsMA/wQx89TSROZh1HWtOVDh+iw/purf0qQH2f/lyQVf6ztGF82JBN10wu1qR0y
z4eQxkMzEY7PQJaj+ryTy4jug4EyYq04pRrsdRMO1/yev+CwcqXODktsPBzoaKnD
ujjJ8/KGgIx6qO+oBY9fxX2dGAgF9dG4k5Ahe7ehzysTtN0mhLr+FXm2blcuCZP0
hzyq2Ue2mpaWPOQdCK30xNNP7IbXTTKSdRWzn2R8DaPkIEJWOfhy0D+huELIvHpG
lttcuu6jXV9T2RWHmJ7mHHhdYxs0Gg1/yVC4UeI7brxVA5bQUbkisfvz9wIC5MB6
ZAOYnirKVEKcwZmFGOJDPhy5apEGqrG9hJl0rDSQAa67uCzylcQHXPDKfV16YzSd
9x30bo1I3GX5OZZL/BHMopSgN6eqERDI71TBzfEbVIUeL8DpzTVeDTiXWlS0yqer
k6blX8KEdvCkD8oEGgiZnC2L85qT7xi2XnDK3CH0b4nhvLX0xveenICTcnNwTyHJ
4bMeS4hPaNODeciRizs8LKfhRSDMRKAxTgaqfRlRr9PqiIHJxxjACXaFErfS1iL/
5htVtB3W4e2ckll8JFrFBKNbtyG5oHz7OK7J2yh2Ve7Frz0pagmiSv3GYOp3xhJi
VbDetw2no6KrGGdkXCWAjiir/RPAI2yanCLVkghEcexWqSJIhNCp6IdmRirYSKg2
YLtWYdEp5gXpLj+y6Mn1tzbQR6EzH2LrUuWWX0KZ8F/CS3zRnxWRDPrlW2MIG+qH
d0JIX1z+AE/ZvwOd5/Ke/xrcOy94SoYYDETWrI1wj2Nf3+PAKz4yk/eh5/TVdN85
/bBvtr3FCCSGvVRy55fVoAGwo+ghCXjcAX0+89JywsLjJ2LMEJIvlJ+QQd7baG5A
SXJo2PQsYNLa0KYVxVsxyPs3hTtqKvkimjkjzEaLa534m0g1gUG9CZKykb6K8S/k
9V4av9XKafpgxs9IxLbKn5ieh6kQ8OXNtUi12gdd7ZI5nM2JD0G/ZuoSxgrc+dgz
bYxveTBby5bAsa698IkUKQ41HJrIw3SjoiHjTXvaCNs4CdWhinngvCAmWztG3UCp
iA2E4GhdlGOx+pGCBadx5j4spHZOA4xZINUj932ZpOuUCJbbQdd/2Eraqi6Jxdad
vU8vuGYeD3wsbgiczwOKQ1qQCQOdD2P15pDSf6oHYh04+U3HnWHawQ5uvj7GNvU2
LF1jgDDNHidahulNrIHRasGTUFSNek3F4znq2bq9uG+9LRYhYe+mNFlWnTf52JG2
UyBGYcouZ2QSo39nBnCVbEJzAGlthlwhVJEBjVQREbfbbzPGKxlckRqPqSiYyNJ+
qlbmEb3xEJZMYVwVVAI3tj8P0hNl9D+ctXk5IfvmuNBslRGErQ26WyNeOT6x9VSi
pavxT85nacOB7fJDTd2tKbmkQpLvgK0q0dw7Ls4E/6BsA6aSqdXZaJngE6MlX+3g
XqQNCM+MnsbFBth/Jdol3Eu97/qhW+K4JWH3ye+hrLvZcTjoGtNYKS1HfwGhAV+S
csf/lp/WrU7llrlAXxg9v9/eW8reuou8i6a4rjBpW0fzUq5RGjoghazfZmF7BjbC
WIJxhVIpBC8XhJG9TmNQa00fJJD78MXsm10y1TZW9lGRO9KrqpgEwulcZdRcjRbL
Dp/LCJkER/y/nTYclBhbUvxCilytTOAxtO1hOfR0A+pwrEpX4OWh0IjNLWBX9/Tn
azGXOTShGUjv+5pXiIH1yLllMMMEqRiAaZiJwczYpvQ93ivR8b81+ikd9ymPNgDI
bt5c+XsqoxD9UPj2kNbsILdjOpSmW1VkEirUp2wEba7YChf4YqllhF5elQ0F1SQd
sLdl2LA562hig6zV5HMBsy6/3rHA6DY3gQ3kKRz+Mm0Dghe2s9CEmJniDOo1JTc+
4OZarSt0gIKEbZY+51wCsW57hNawSm6SzWbcfTBZKaLVFA31d8XiqDjW1Yd6lef6
DB1RrJ5dlYIsVydXu+9KYSG17Z4ElABARy5rIbV9AJabY4tzkh5/yfwsCR6FDjaA
bzVDj5Tu8yUfbJxvQheGLyLuT2U0PlBSPkwCbXvR13hKhqXNEyVN2UkkNVzEENBq
kFmmWBgwIyvX2wWs2hJUp/u24rtqwVb2mayXRC/X3noEnBOvICn4nZOfngOZqnS4
YekWtHKJbSi2r0Pr5VyU14dIhMDG5p2NNYkfZ0Tzruu17lrRB22aYI0lPUh5fMKu
zK3GCRMWj6HPFlkUKVoj2hQDLMhZdvVOMOQYJhy667RvtEpQppBaeIcxXroEmJ7f
+XqRwaeThkfQo0CmJuuZmTBWYuSSS3l4KNn8mWVHlNKM+UMeRnJxcXloxskRQOFc
umK86tyGZpvU8mcEdLID83y2LrNkl3QCdKaR+SITnbbmvmxfw94bjIgmvnjjrwZA
8J1JDySX23CwnFfMwnlwuz54mqXZA3158vCSvgCQxRlF5iNmEvdmLx5mrgtsVswx
4k0uEgYyuXHaWiEtj7feuaozorCxF4iJi+h9TdKZCoW0fm9AnjYjJyEudrA5vzEz
dlNCHxGWf7kGQB9sQVBaIFkUWZPEoSQfzDiLa4lslz9Ua16kyFvJfO6K7jTkK5EY
DHcP7ziJr6m3RPv1k4xur6vHxl9QF1BKUBhoDWdK4w+kaqPctnfe8LVigH8jpHpm
e/ui2ROd7Ro4pzK8H5exR3rf8YbovQdFr7u4WmpNyQnTzMePV3g7Bt8Miz4/1Owk
9lYbklOuUwT9SC20QrAQ/AYjuy1wVPupBOmYZvz7uIGT+54K8ukl/un94OIEW5gK
atkKjT7BrRmyXdVY4jaYo/yAM6VyPNs8pTVo04fpxV5rlGOcor8PoKJujdasxXtL
HSJBFOcQTTrmke+5Q4ESQ14i2Maw4RQkAkzxy6rPhDnJGln993ve1TUDj9NM0DXm
Luf6w7KFml3SEN3uwKBmwTdWXOMzJ8bpcPSpXHqZ6uNDePuSESteksHgMU4Mm60q
DmcunTOjtfvarquXeIQpsRS3b2en18FnIkvi6BXhUevS6jrU6G8RH8josv5FkIvG
gwEmuS4GYXabJFp/xMyQgTNUsYv2gcG8VtltuGKKgljR+T+wuSIGX8LLGaZgQwqb
8FB4acxP+F07zfliJ9t7wL+rOLS9avlKvd0g54MKwLqSBnJb1/2YIcsSOcgeTyIE
2Nl/Cp2Y7EWtIETp9sXkCYDtpCk3VV1S51YnW+Wbeh8nbSuT5Wd2z6dAbJoCfQ1r
CU7G0zqbvg3eY+pTEUMjuKkUR+ElEXSPeb+xILzQJ3Gp15ClgkV03eNCMoRVgNZR
rLthAk9tOo3tPBAdBHDazkOUEne3dFmvu+fRlySJQQtdFJa5T2qBDI6JVSq2nYQd
OQXurHyLD1VDqEgeBbXr2fB5ZKLZy7QlN1goQSDFQ4DszVw0LHmSyq/Pkn8+XXPl
hXDkEy8mtgpzT3ZqZLYu24cg2Gqyq0IHWZpSx2RjdtjaMmbvnWLAUtRqWowmxZmu
+VrqS91fZwPBZ//+wzKAX3JLHxIabFI2TF56Lz7M8zWFVfEY/BxD9svsy++E7kqx
mQoXQBBaV2AMee6/KnD1FnPHFq6E8SOWByM83UHAH3FvsFXtjFOvBydFZ2YlRom6
bmH/24qChwecw7e4lVyS/BLmkl+gk3nD+rcNtIVeNN4jnaCnshVlsgFOO28FtFrV
hAQtu5QWPDu1Pw3MrkOTR+itn5+NNJyZ9ZfOcqK8DFNRqoiFm4DYIdm7E7NiTlX7
2sc7NpnLdPwCeywiYErNwyQ+GyNE3/znpODww/50UG1ilb0Z/uIafDU2UDtu+/E1
waATuLepOxN+N40HdT4NxAE3tHe50OIFwxQslAA67UwGYngORbus9Le3EYhBBFng
efMUS6bLaIg8iNyR16kRqHpPMj8UYG2hzWPwI/VFR4CkSu8+lq93QTamWJRZ6wKC
21JO+z7/v60+5Ae4D5Esz5Q8ngbF9Dy9sw8CxoTJBDhaHu7z9EKQ0Gy92qMtqKjI
5OxwiEQPcl8EW6HHVkzw7F//XeSk0GDK4VAePTxO9HANrOQVFmlMPRY+ALB4NWYf
515tuSQDIrEKhUJzqj2nJcZGwz47tKKBBXyHirLIG3UoTewS3KaFzNbEyMKlSJFe
dqHDdhtGNFkJ+b0U8lGggKVAcl26f2Svwyv1loVqrHP6BEw3lEMIOvPnsEQLjiGz
TSZ+zvXvI5fr4pLGgEb06M/uxIv2FgzyCx86cUlj7Ec61F4R7OmaI/YmPzCI4ZTg
MlowvSDTzfn8sPlGZ8xAevF3xFCVRW7F6g/ukoCot/zRYCSqIMH+WN+VLNIhnIml
p8C6LRpp8rT9N/uBJRUd/E99+hegMSySrJiLepeUPQzqQ7+3QP3CRWvjhHyKMTBs
bhI7abqpTQOn3/vBnL+7Zy8OijU1sG4qbD/PIbbT32po5TETc1/951G+GILv1y7J
tVNPfnPJEuu13FeMh4WXWBysi53c8iNK1B4/Km2vToi7uwjNaB9Kb2cKHJAuE/qF
ZarDyUwK+wt2M6L2Av1WUAtuX7tFDpZLp9xHk3lvnLc4BpF3TBDHUlPFXog0b7XH
Lkg+O3EED+RSmpzuMswuS9UMsj1et2JO/9xU7oZc2Aj+33Yt/XHMDy6mBpF9uy67
M6bRUuwj3lEyb8zeSIWyIKAum1MqZNU5xPvL7jIqKQUel8A1FMFDKSr4qyqDGVK9
1HPSIA5xyuzrdZekCyvC7czzN1JcutQlsDrkz+8hsemUI7muflfjFSTNP2JNxyiW
3418hvWvsWm/hkRKzAcwu9tMyLdKfBQtnQtIvV3zoBy/jGKr6BIngtq2kTcZquZh
GwjbDQBNWAeWkFa4hTHMSqz6Nh46gENJGsdXsQNUp0cqko6AE1aFZqy/enMTr8un
ANOAVRIs53Dmgnp+kVUARbw6oWLEropyKRtntBsXDthOcbvmX6jNDBVk+4Fr+sgA
s1K/p6qLjtFI3X0uRKW+FXar5gJ2yZ9cwd4zZ6IuVzWifpnxNWu4r8HKVQyU91r0
WMSyHu9v/ePWbuHzvc2rYBWgQdL/Ton/Su28xyVllukILj0LxO+2Pn+0iLh8pzng
NtOm+KOiuTbmjYpHWEqiXROiomUQi34HWTgmnH+CIuDkRjDw7bOut2C8E7C4skF7
J6XBNwlGvnOqQIWxlxRYFgLcGLBuPvoOOeMhFvfS5m37b2CFXLthTA5ctSV+j7Ks
fFLd6iETLXPoG8rrD34crOXBdxhgn7c9eQcKVN67YKnqbJDX/nUNHN2CiBUrQVDt
033oeSHfAVQqXwOx6qb8Iw2bL9zHiNq7wcAxZoFZF/I/I0DDNQNAfCCZxY+aHLMt
m1MdJpUTYX6csXonp0nqTPTu4xGT9codV4oC9HMbQMhA03+yIDkp/0fCi0cE+/g1
YfmZ1x1IO7Oz2kw5CGJ0qzCfm9jsriUaEJTqcaQ0TWkJcZehWJRu3G4cduIP5pzI
zu1FRt+WlshW7B8pdGye92l0WvMstSeJgjrLwTtAF4gM0qAbyeoIc5dJg8A260xX
cFyhiOMC8YphE2UOsxbzKQ==
`pragma protect end_protected
