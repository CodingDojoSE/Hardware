// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 10:40:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Li6Wm38+HrwqjFxCrbaI7bBITFOdu+4o8DswdlP3mZsw8uHakY9vf4585DJlO1ij
PpOqnsC68BFjFpAUOoDNdddZ+3Hjjo8l6uHTP8ieDjtTh+btz9j/H5y1/256KH2T
RYp+T7pmCsc5hsurVc9xZemCZ4XBka7WIPQAp1kVaVQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27920)
rrB0TavqpQxNU3nBN0oz82/PkRn0ioIWtXOUHMD2PGqFM1zeQq+DV9jR40N2SPjd
0xbkVb03/Okb4gNhkQobZnrDTOeFucgjbZuACD0w3SkIAsYVaFWlSUlpxf1y4H0G
urgAXGPVZomNPphHZrHHAIWA6Eucp/mFeTMa3K9qCLLVQ9lGdz30rJVpBIpIlygT
5oVRAOWDRXzWPXXRe2aTpqT8M+DX39LL4z/tAdz6IM3GD0sUsuvfHBYyfJAy0is1
6avBHqXhpVe/QbuGa8jOMc5WsOhcDK/28O0bj3DLw5rdXlfkLfJOcrpOQHXpYkT0
tR6EjFHeP/P42b1rqhWIp/ajkR/v4tZBBQXrZnbkZsZJVxDJ9YCoz8BkBDTbQieU
LSeTDTDy5u7Gd/zJNcpR2q1mdajJR+Y8ENkUyDjnmS1rskt4AKJtc4o69cx1uUvm
rXL5AUTtx34pw9A1oW+K253juea6npBH6L3kvmzpR741DcWtck3fDN7M6XdyQfWT
tRoQe+Vv4I1woIl7wn1pfVRnDTYUABiFDpCG2AYYVWd+gjOc7SNNcIbBIsamKSDV
Gs39GYzXpA0s9zH+gK7Y72qs5TSXKhXVBoTyirKhuVlTqrDfQwQFvoSUJ+orpBVE
W54mvsmRi6xD3aDOyfOAPJz09YXF0QABh1wxBYVs4WnB4Rn0we1A5JTNWr8Sb5OP
Pj9EC5jhNBauhAISRfmldWo0m6BHnJdQlN9dH+DpZunb8eycoXjsAVPfbjal7eSh
HNyc6p1i+xCYjo4CK/MhLl0kfr6wysu9jgH3Lcn/BGNoMWwlSCf+8zYu/OnoH31I
Jh6+CUym8eMzskGbzgzm1n/1p08z0KPQvJsYhDPbsCc8AXSD+pv4AF3DzdhffrZw
EgisZyvRsfAeV88WhAAcbX3L+ZdRFkAUcXHGmQ+ttS+5tar2HpQyudw6E2kwUSqu
AC+uNP3nmu/sevSMCaUNvQcpdnpDubW/IshX5MGSjn8t5wYKnyj/hrTXoAKqi4De
oOeCqfmm49LPFhzQK6mfPAVJFilWEQsRPEQqQutwyYQTq9PfKFnCVyisZcYj99u7
3SBLU836y1exie47nvTV4ih+pXbJGqITbUba5F/J+4tVfpwYgcQLE64w6HEX1hFk
CnNsIBRyGe++YPLWzsXiIDpbr+CnLjqtxJJtDcK1uKzyronqwSPbz39mpQUvUMV5
+qtsBWghH2G+pW8KNxmbPyhLyLjrHz7EEv+sHq0ytQdkrHtAoqx0HZQak8Ip5l7x
WL+J1JK/BvYo1zrwMHohfpXfRXB0M07HbIc6lJwyO402L7Mxt8bJGRBuWN3ZH/vB
6SwMIjVxVbOPzRbu0Ez3ycriYJcFyRpmZzffBtGI/3/2sB+MVZdpgCkF7f8WkBP9
gyqezDRJAzHlJ/Q+AGzNfJRbgnqLHOqb2lYljYqM21W6sQT3mbqnWdwsSMmznSYm
nXKPx2PCCxUcGEPuz9Z6zCTMr7dUhYHGxoRg9jrZpYWLRHt0OH+VOTuo/Q1F0mF4
oB9sK5dWqf4LQlplMT8sGeFRfWZ5tbFaF+JYuAB9ykIIiPelw3R3nbKP4GHbrBnc
iHVJUsN7b363XDQ4Oxr4dpkpYOLFUmQZ/Nbe4DJETbFEJjBycxmEkOPT2dwp3Cij
kK8B9nO/C644XU9Ec85yMXu4mMResJnC4f9nTKKy4W0QYdlpuCSVO2gub6u6YjPd
eruBDFgskig9YCQbF5jmvCBERX7U9vr8bcA+OH+Ruk4Q+jZs3io9GWIdN7fcnv8b
ADdiYXQVz+KiVeammnZ9TguKBPMcMjAu+zoNyy/zkXBMvtY1Ae4/4hlqAImgRrQ9
ht7dLNHnu06t14Jkp+ne/pSFc242asOzKV3Dkb/Fn1h2fsNzulCK5pwbjCzFcCg2
hFyQo4ybSpZbDp9ZwX3COWVzkpioZDDL2NQeaUEYm3vAWuauikxG1v4QkrwZPxcA
8Cv/s6jxuWPWC7G/aGBLHnHqmkGgt0ran6n9fj9bYAGFWjxQW/yeconP7lNiy1UY
mg19VASOosUIUNvhSNjQApayJ8PBC2JkWwlRys2lKADsbGOfdWZaQmejS2qCMDwq
aEce7Akx72zYjnm0Y2kp/VRWlrNTr1GNFd5MkCYCEgMgnEwf/O+DRpW2qBWDBye1
a8NFqW1UStcfvxqUdvYcdiV2G1YD/DsEQZoG1jxTSyjoEZdQr4Jm/uWEzD2ugO2Z
Ylx701NAEfv+sGSlBIj02Zk9PAFgZxDyW3mHj+DlJ5HpgqPBRRhcaCX2uU0Ui/X8
sSiwUQVXAYM1U02dLj+x8E19gC3WOxink16ftKPJyRPyJ6HWqTAdvhrvONYd2Rcn
5qG5JtWKiiIqMWFmPB8NluyNXNWd0ZAAL+TJ3rShzIAV1sN/8kQOxeqAPFKG3H74
JYl9lx7UZR6mXnVNLri04sBAKR0C39vm+SYhpk3qDlEM9jzzZfkRRtZho8k2Roy1
Dtt9xrDokxRw9DqR/R+VmKfXug63srt30HlMd3TJSZ18li+YBuKBiuG0S6PPFC7E
v3Mf+Yk+GanqrD03jRMxLJNzhFSaKI+aYYN7ZTO5fmwWZD30bL4snGCn9lJuuIBA
L1zfY0l4iClIItOcH01okgg1nsZzYk9HACeI3crYwcZSbHKBE20CGMpnSBA1KLTJ
XxCJU97+GdtZ/hnD1HZ7xJLFQW3EKT41/ZLBOel6BqFauNieJOPn+bE63sW8loBk
epNgSk4FnSNZ6e7nCTH/8pgdBGTNLMfZl8JhcdJdE9R1NJBH+Fk2PMgqgSbkwSO5
Eo0+VTBXCqGVrRPx/hlCrZv1nEQ8nYFpZAmU8TV4JUxxg3szD4rwcZLQVUZXxQ1u
OcTgIuhfHFEI9wzUW1UE760TqbUfQXiUUX0m4vHewharOpOBXPxARLnMwzGRCcM+
hRDorPYDCAqLqm00TL/FrT/A596lHvyixX0KmOSFv6EKL8J3uzRwcJGLZC1JqL+7
bPpJjvWvoWqlxAfZS9a1+faYU1s210YV6AIhMMC0IVjglKFhPtXdxu7xwGNMZQEj
ojqedsITvTkJqTjwNNyNjaBqW0fIHlGmKawMGHjJV8AOvtfwQzetEJY8aSe/Wnfb
05QFoDbFolD7+LJn4Zm5bf1b5RD2Mqf7rAJeYbp89zXyBlvDjfu2balPWX+NU/Oh
5GSEtZxgx2YMSG14jSUtruhdtse0EWlDLRVC/HDT+q03115EBrX0OHQkjtfDX+77
FhO8gSSCM7+gYWnP2OghgtB2+6gT3RfD0Ean/5tHWQwXP733GAMKQVgfNLMEsEI/
Z6l/nZGnllwHAfnR+I3l1Hz8Mqj4B5rywGHW3mXS0BJqKwgAaOd6jmuuCcyRGbrm
B6LBWB5e3OZ3xXt2bIBNs87KxhJFKEWG8g4y6TzmSpasYp5tIGyyQyeqScL1kEl7
wb9V82QzQqs6Ub5XC5ZPIG10VlGJA9tXOq1hgF1qTUVoIP2zNoWyIKdRAZ9nKhQX
cLsSDY+y+xT6HzrL2kRneeHxbIHWDR7ZekZ0VL45e1Jg/g5kNc4iLYc/ZVUSzP0O
xgR87YIcg3ndSCYVUpO1EZXDO0ajjQA37Wzhkp31wsUfEY6oMlqWJzsKGx+y6Q8g
kOqdNCF7PLHMkG9seJfmeP9wAgrJhEnQWOUNjqnH2/MWCobjkRX3pqSJNGxTkgdz
ECyZvzFmLZ7JEUdSrN79mUOq/ZVsZsTOFfdbYxZkRGoKgJhDeRUo0IwTH6KRta4v
YDbXlVdf78j7dGWHUFJilybzd6PbnxBLEoAGnuoC9XOQBdaXXucq1h4pZRNSeXGh
eZQn8jGRL0Hi3ty350wdxM2x/o4OrE6JPyk/NTDnQztRcKX6Nsr1tD54i8dvBC2E
pINi+V2otWXn0vwscGQHtyUlniKYBlCoAIHbmkj6jh46NuXoxlkaBsI0fHDeeBrh
9h2yJ1sczRR0U2daxzg1x103bPHaYiG5qi5jHQ748uDu1BGyEQmSHb8ylp+wS0la
ADrwSai8MqXSS1uZGCzsqd5tZ2PWGFPaFJUfLcoEqBufiBKvYG1bhGuXv0Wjs+e+
RfnfYeo8OZvHu9YVzzuaHBXOauF/Ax5cvpHOtICcQlRLqUpSQn+kQ3Cf6hfEcBJp
IYuAgWSSeamEGlxXxwzr+R8NCo5xYCsPU0Pds4FFK/ktyKTThZbtaooIrOXFoZli
qNd5kTU9juzER0JETfT+VT83IzgtwY5cRJ2JjJ7J+VqkQQP7zknNgO63lPKIcuwd
TBiAzFWYUke7h30ZVSJMqrrw3K8R3i0ETOm9es8CpTY+oXwxIpXXo8lg6PnI4Pay
3pBC6C194IM1n76fkNFQr6TJiUEUc+RorSgWMtN5uutZns2TsZDQvLIJ+MGI0Ee5
BgZAdzqYvplcxiThvARKP2wW65oZYaakwV9+YkHbgv/1SJuiQ+gVouDyMwHafVCU
9R23/3Efe8JQei30lIBR5FWPoWnZ5iz0vX5edh7ATKLAr93k9n/4V5gKs8haYZ9/
As3F2S8e2RJzKRHL6fvsTnWtMX38ZYzMiUtGa6kZZs+Uw6Adcs+oEkd/tUo62N61
FaQkxu5rMBhRtMnyXDgOT1LAURE1MMQ4Z3uJLw3r3aIKIV7rJZ/C2hyBEdQrpNBO
ZzYM+nG1qELhEa5pgkOXMt+0ECNBwgHjrSYjT2Ou2Y8yYotsIBOwrlGbu/6+BVEw
lSaLH95xWFoJuRA7cB7f6VaP+958bzkmW334Z7smUWE2pr0XwpUdI7MJoW64X0bD
KkkutTnEPCPE2FU4J/EIClecldo4rIBecHcsHDr7ac3fOPtu+BpN1QshiaBR+tvB
vsPOmITYsjDBNSnGxhP/KOrRochswhGB/dpyy6rNHRE4HhilVzOMnbbFj63YEbN8
zLfLGHzH+/t23Vl49G8ws2Ys+uoe1swYmeSOWH1oTC3RGoxWPOa9wUidP8c6ZaYU
acDu1Oca5AMYeR1/bEr9CpFQ6qhQVNKAYmVrSSIXTGlDd/8QKfQr/HG0F7LGbStt
GglwAsaE1ksz+8bsoEE6aWvqydlZK697nmQct9JgNEu1rvV73rGTjSSGu/IUIaBw
Id1aL6hZjo427dYU+zKIZMkZkFCTtGNAglf4g3UHDObQYj+myJPKdGcx/yrGEOmy
q16eESfdIQPMxo7u+epSt7fCxVQZRQZJnQacMZCkDBxpHqIfGVaRdyLIP1/xrygz
efkHD8mFgT38ULGshe3s+QCVw56NFf47zGXgpYzONIxfGOs1M+RETvsiEbGA4TwH
7hR9oOQjs7szR2o5moFvmIWE4uam9rSHDSIflWwxGl3nMo5E1A8KizdQucUFTlvw
0tIeA+SwK9tEvXxOCL4eS00dclKRWWgkWw2gkwwz66Qc66B3KT2oT6hLB+yjoX9N
S4rI3zU9AJLslJA/utppfqCPPK9GUBJL1uuzyEfFrEVK5lfI0HKll4vw8TvggCUN
NkTSD4CeFWkNU4muA+v5gY5DncX1prWCKBfS/IiJMF6FveFgU2Z28sBta5RV9lJt
WBCcIBG3Njjtg1Qr1GlsS7R/KvLtg0ZzeCTOzdkakciG1ezyJuX79PQk9s/Y8um6
flbH8CUhb3VgGbfSlqLLbMBM/GkL/Ixv4pWf+Myei4K/PHid8TBOrhB6RPhTwAUl
w4wL0Qd0MBQEucvSnYQ96mT3/8VGv4u/4nhCeQEulspWPb58xLcfqIeBmh0LrzE8
GsdytUH7QefxfdNQgufPvt7rRBPB+phNv8C2Z9z+xQ8mM51nLRldxLnTQP8fYxub
iJxp3VQBLJLIjL1FkXCWVokr7rgHLezSxuZHz9/EO18QSDyQ6zD/rUuGPBdcudQq
SLe+BSWd8yssOZbUsECxmm0nShqdfzLIVJIM5hw2YT1CzlqaLMPadDnRhD5jJYcP
DwNGjVFq/AJKUE0CpsUcmMDAykXvyWsWmb0a/8BopI+0iw1iv9EwI8ImyR+rKQ0t
u+wZBiRNM/UXTsJpPGO6eAz9joYyNvZNdEeDskv84ot1qWqERK3HYAgQW+tLwqXG
YTPdY3CtHQY/O10asrZcAM6QZP8CYGN5OxorldBHkOc31lc1ozADpDszj95DPUnX
oGgOpXMm5cRuoSJXmSxCfjK+Gw0rZhquSk04kZsAWF138LNYAVsIZSiTRcDNR5jD
29BjG7hKZoN+7eYMwtUnoiTmV60FL7T6k8tZ5YR9ILAwioXr10hrd/akOhhbBfAu
UvmNN4+1j7D5R+NCU4lmEQPJyCPqRq4IL6FEGbun86fW0ijHLvH33P3HrljLBYDm
FQnn7GnPBJ/l8cqPm2raiE4zHJD0OzAPtSywNU7So7eh/+UZJVWq5HCyA+cFLkX/
4MVqs/bM9bl+4YxYf55bKlBfQyOHxc6+cHgNxu1EUaReFedvDB5WPlv026Lkw9LV
ZIeANpuJCSkofH0+M9iKke7gLKJSqXq86fkXDeleYMdjQZY4glCZxUcBaA2wh70M
QpT21n4JWc7p2u61X7h9kedZ9N+16u3hXy6/yjOjr6d6e8u/LlHtbTX8VWUvJ9z6
l4QdevziKBH+cIkNlqxO7o6xkMaoXl0s+tm7mbIZ/NQUoXUbDAVAOKdEyMOeYOXw
0as7N+gjNKr0yIeH498zpEK59q4i2EpNtu9v5OTb8IFeY41RY28aC039rgdbQab2
T2wcmcnjtHXF6xTFGGUvuyAFhjXjH7myLcqfey7PJhj/xj/jiF5n9Gtk0A6E6LWI
VeyqWcu0yBk5zJf8Ialc6z+SgPe9trVlgm5DBvHPi4OfiQHmnA48fDH3as1zrnfx
VAc3AJ89fFzmGf7sE3VjB3zVYqD1T1YRn6vKEs1mcjgPAXMVx/WkYEtLOnIh+isI
Hb8Iiz3AknyeKEcORr2zHeQyLfqdcGAb+3hiRoqZE13KASHkt32ks7NOmLx6N8vA
BHUSyN/n8KaXsr3oYKMiwod4VyGB3Fx2sRo14fjmskmIasZmsg4kvcRYXlJeOi8/
orqXtN/ga1Rdxx14rKxRqcgPjBk7yDtuBV6wD17zdD0CD+deF3hIYqLUVskDj/0N
PLDukArztKMGQ4dvfC7FhKdPaeeelD9UuAi5kL/kgVpqo8mbqS+hjz2yFh/RPcRn
cy42M8wpBBZx0y5XHhdRxl1HZYiTUcy+nZt+iUY076mvLlXxgwc1RWi/iLHThYC1
EW4qUmsetYOBiokfY6PbEgr4RkbQcGOzDwAPK47RhN/sM/kcZEOqBuxOH23IkQ3J
3C/wU5lfTpJRqk2BwI9314GuYankqi5/yi38bK0bpehOOBghlqVf7u3gGU9A1e8T
9IgFN+SOOp1HwMEdoa/EnOayDlb8oPYVRSckoFZPTcCFPmFpyxOaPJDhQHyY7az4
Q2gbthsS/ie9gIHHAiiv5O6kyEXp8Ec3OWnWlia/is7uxBSyuQhrsPU6rPZw3/hn
JHBAcPOECanBpYAd4NFevuTlE2DzE2TXzIt9OtUvKqoM07g87cWVFtLgZuevVLRL
kFz3DpBloRyzhhj12FkLMLqrF4s8QshRy9dwp6xxdZQsTcn76738dIszbuu7cEIG
yMH8TneBqvj8f4WYzcHUtcqylWvYcBSA2hVbjRS4kFBccqykttodFGnodTmD4Ida
mp5ZWtRFWy7u7sp+ulFzZluepn3pzmhvMEfSVNOFGVT9Ofss4rySe8Vr33WVq97k
vvEodJj2781FIOKdISA71cSXNuOyeDrvitdUlJVckCEMnghKewlitAtazyIWk0kZ
+k855LdPPWDqFiQkyz3uq4he3+cdeX5Kmtzcg0M0nMnGpiyw3VqRMwY8X03lTAA4
K58AMFXtKMDw4ytLBd7ks33UibI9UHaT5g5JzICGJ4aRltHVCo49NWO32rLCir64
v/W3WHqQp7hlYVxWnNCdoEZC42kcl9PE/f4701p+RuFEbozLLW3BBJ2PoLARTUkA
8W7Gb4Lo6PIqpvfDA++QgEFljcAcgu2/qPJUAzSyQDQgKretXKZW9ggDdWUSiJ6C
FfeaOSxs2Y05wHLWbmTQNiB5/nkzbLww2DANXA57rFYkediziIk/L/QBXrDbeuxe
VcMKRFAJPuJ0mG8NO/+1bxF7gdGhnRwLP23F3q6qyJ9yScsj45r4YDKAgGOTkfho
j7GgYkhoKT5THmxFS1by9OfSfi7mPewH88l1Ul799IeMZeHBUJ1Kcw67mB4fZcJL
7BCkHpPM1ZV69SGVmaLafv467pTAvJsdDerN5EIeFF4LsdiUecW7Wadhv1UtAPgW
y7342ie7y4FegeZd2WXlfect11VjXn2YE/vkamGZPXUmYVFBreI1phXH2DsEHx7n
fG/n5mwYKUP0/ATZhDzJ2HjjUjOgXrdyTkP61FMxVzGI4vmu2Kh6PTwzIKPh/s6u
tOHH5m+ULP8Dca58DpieyfjMpXRDk1nDBBQzl4cQO3PSUtgYDJeYNwpj1XKE5/RH
bX4/vl+8wDmZA0eZH5GnTocBDNnxgAjPzCd10NtZJ2avzzHVQMpEY7nVX9sYpUN2
o/W2S5lcafugJAYhY+SUSn+mNAgFKR+fXDkI5IMdOwv6GGt4uMCpLprnuNHkDRtH
ZFQLuwOAQ0JPIy2wqcjM777KUcUfvOOf7OP6GJ22uRC6dZ/Dv4cl7ujPF5dIO84s
vYNG2QaLW/RY/6WMle8tf67DN+/7BgVKh/4GW48WHNwGchJHZ5Rzhtzvpkb3cpCK
J2DZOt36EhG7gBs4i22XVwtSwoeBaOZWKWKyrtZGImMPknQy/YSRsNtLtldIyv2w
uxFjLoUFCzN7OMgre6jEWPmm8JZsMxuNCm8CzGn07a9x8YqhCDn+LIBsbjxj3KiI
oX0VSpMmdAZTQMC5XzdhlmKZKmdiEc9UKE+RN/LHI2hWNhD7lqKZrlZJBjwOvhug
Hk1X+bybL2N8drn0zZbGYLm1IhnG/KTzMWGrIQsz63YdLXpAPZhF8t9JhKNLGtXq
p0/Ba8lEc2acFemJWcg8xjWgglLR+pnXs8K465s62wyF1KSv0wNJsGhyRiv6i77b
SQtza1/Jl5PHvnLC4NRLAGC64oZ95UdNb0O0L21BQIQCOF3nhyEID6xJkWhbB+wl
S4O+MDjSAJBOguWrHGRYjAdET10hIT7aOQxHemXjeBk7wP+aKuTLxg1USgjh3TRK
3nZVlqgaD+rTzddz2NBfa82CIrw6RB4Qj6ysA2Md8QOZVO/ApOHBmprR84lWr9DG
co0TRR7W4xV/WVhauAiHRvN4dic3i4x4x9WnRS9lcM6Bo4ZZ0TRFK/Gpc/fzzk51
Oev+o80HkNoWBPZRYXiHeFrXIUUqKAIiPpJ6woxafPR5oaPtC33lMlcToZzmd3lM
+gc28ybJmA7roAuzsXtwVg3nHMG61nTOViG9uaT8SMeq7mBxvUy0nTpZOMi7bItA
kviNAtTHg+LP0ZRGT8Kor2w8moy90WqFHT+gtGLn+L4Ilx/dN1pKQ7S7TGx9+/DR
dapO/5b+vH7Tt17gB6fSNNtUZj/ctZvAHGV7RB9QfDQLVjEVaR/TpZaxs72pfcWo
YNWxW2A9rTuywGybIgd2ghCoaBDMi/qxmjmlsHRnok5i3kInREWQQmI38ZkHkx/A
EwQZRE73f6Ehf0A/ku6gMUTqvm4dDm6a57pLj1EJSN06J04s0LHzypeVWCHw9doH
2Z4bumT390MCJLPlY2fOH20eC4juq+JeDImTZ+MZ0+BU9RC/479t04uHJFz7NuEO
fofxBmKT8RNIrKC3+Vr9jEH3dat4fSI3zcuRQrZCVSO9DYuEG6XS3ifE/2quWIWM
FYngD+czEbueY+uDXHra5/uBzGoWpVUuME7w2q2NK1yKhWmFd7XtabsWg2/6K1s8
in7exRrV1RtQ2gxrShhaB+c9lQibwtwzATkC17lx1az3ndSYZ0PsGjQr5fuNW8uV
1K/tWt9Xgg3vQueBmwLWCYovI14DR+CCKkxo/AJE5unobXt/bVI6C1I7v7qdWTz3
cmljQa57Rff9yJE58XiDXvMN6u5vA1qH2P0aO2CUsqLUob7/EliKT2uZkJ4OpgSX
ZxKO6BspDRzX5YvkBELfa7X3GVfBVGTECVbgfvZVNG+H43bQreAECEniWsgs9mpC
n5TP9GDb0l98y77tkufhLtIUokUoVYZcvp1lXBy+fuKLJjWj5vrRW0MuE+t++lr/
LuFHQmabqovmStWUJVC8O2QC8mM6H6DFVst4gmFRrGJNUO0JV0ezLxjgP4Gi01ba
yh5A3Cu5e1Ij5wPqLiTsmTaC2F2amxR3ucFDpFQC5nvAcIdgkyG4R98shhm8+2EU
q64IAduz2z+y7VnrX41P1I9daPuz5JheVh5BZRUZJmZhhC1DX8SsDkZTMoWWbh51
xtJa3MzT0Zq3qyNLShOGd//AN89+6F0wZkm62hbJNXSFO4wBmEwX0HCFM60PH+3+
tE24gWcBpDSSU+d72Loe6x4AuonjD/woZvCIclvhx3GVwE4CpgXi+tbBvtvf9SjL
074Ggz0FKoJOcO1xOoCkFN+qsgtc65XWALBgM027i98yxsnpGRIpuiZ0BqhsDGjo
6ZbsS8uRyfduGblrbKnfvYE/qXC0CB6QnoXaCBFnVmPGc4NCp46gZCSkRQSXdL4M
0nAiCOy24ujLn1xzqufDxefNTTsfy5Yyw2Sk78kY1p5kyhkjK+S+IgrAzvDp8M5O
EHwIqCPU7/tBtRn5hG0UbfL01Xvgqyi4cIWKXHgX6wX5p6A+LNusHfGbvfxtdyD9
d71fNn8pZcblFRIrx3UIhM0kYp6WkIG4LyeLXTvNIZlaiG7cGbWUdL8S8Gt9hMoD
BLsHwZsdTtbiSKbr2S/jtblfGocQ4OfZjKaXXpmtzDQVTd9mdkgc+0zYpurPQqHL
qzbGchK42HMz+B0XJEonkYtQdENoQKrTrxKl2gF/T/cIqi6MeK36d4+retu53LaE
DNaW12lIy0PeGvS9x/tmzB165xdKlVZgkTdRQYCT1sa1/d2vfD//xnSI+HGG4RDK
m4+yWRydm4jSA/d0Dc3xSclb9UrkRs/THWVWPAUtOoP8ktsO5zoul4EP4TAm/lh7
6/xVLAsywJBz0p/HIGQkPODYTLrxcUqlQ63x28DQWRn0lXeau5oJb9YMcItp48r0
IjK0i1Dh23PmX2YxaAMplBJATrlqyapJFH0U3R5kcvxb1Ip9lNX8B7lRcGQ6ufPv
dyr4rfyhZ7BOoWdZWSY8Hab+0+LOxR8cLl0asGBCHrj2L99Et75lStH0ebgI3sBU
lRgtow+a3sX+UdEe+EVcluRnZ/6Xt7hAPkprKO9y6cMwsmwYx+c6Ooi85UAO3ESL
n7jT3K3AxFk4IWwZnUyg0U4pzCsZqUd8zFbtVnvxiMftmuZZWq2bt5svGtuCS4fX
XTE7kgZyHabXbCxojMuo+uQmuMoflo999R4jaQ2H7Cxth4zIQdeHGfOB6MNVrPE8
Oa+2EQRKWf32OzThozVDHo+o8GWh2P8Hyncn34eel+E0a2RNh+GG0VXiajH9AC1u
z9+yj+9yUaH5xkHYaqWpHDqSPFocyrYJcbRTMztYIBeCi1YSRJEtf2zfi+KyNGY7
VCmliu5KlbTtZv5Ou9ekkICE/Qm8mJ4Be0NqEHVNW1/lJu0unhzZLla/EZF+TzV7
A3Hn5Hxfd0e3FmSbaLiHWAhcjil0s4W5Ri6I6jIBA2/ruLNfh811VDTnwsjVUJOq
RRep4hzT2xhhnMex8epT52TuuHvjecNLx0JBrese53P3CWobVMZdxKrp5Oiq2Gzs
xEmbE3y92TlN+reu2U3yTWHbETg79P3TzsqaZuRx9RNTw6ubElCPoth6nV4MrM4D
ffIIupXqtd2wvIj8dJ9CPCTz+X6VuWH121/vftCSLd8iNkIn6qYF2l480pCskrXA
INYIr56qKw+ZfpHpGwx8A3DjnmqLXNWQ+hYyqC7S0raTL3n5YgTBBzB7E1nxDaMm
kq79QCR82yTSFOy/hBl4T4mrqmHg2HfO6VQb52kRvB8xUaHkhMOenZKZbVihs2qy
iwnw4kgI5CAomCEcmJBUytYzXA8g6ywr3on2NbVBn0PV2EEuZaVgqdIBboW+wJ6m
Z5KN0bGUv8br2RuolU00Peqo5N75LzipX9NNnB0r+4tGuR0HjTA/S2lOB6ZYgaQz
pkQ0ccRiLq2fw/Zg4wVN55pabj0/8f+8+NMTi+JVhvj+wLZwr7fCpRSSUsvlrdLg
kdUIX6ZoziRnCgqog8Zok+CZ9bkDIKvr9uOctdT0TxcqMx84FnT40H58312rr9dw
zz7JANETH+R5aC1++qPe8XJsx5mpHuFE2paZrLb8MN605CSTPuokgUzW3wvnk0+9
uyZta4T8L/Y+/1PwamCglDHVqACZibguAvG6j6iAEwMsm8q7AU8tFzN5e1Lnjna3
QQcx9ylZ1YWqO73/lO6rEupNMhQ3Lo4DT5uxK5WVSYOfEYrfWq8mO5lt8ZReqbQ7
nyrF22djQ/v4pUUJ3z3epSy9l1tWGbZfmq+tI45KJG0+xdkk9Dy+HliPNtjBgJ9g
z1Zl0yydzVatXAurvuqMae0P6KYPU65OrOrIuTSvNX0vB8sqbH5hV60k9sa4VtkF
q32GUhxxugE6zCep+cl/s2lAsZFf4LP8/Yafj1Sctuxk9Bb+UML6Bwj+ulH2/COL
+VxMzkzyZpgTEy+QCkoVnuqfJt6cQBvUd6GDlTV/aFOl/HZThIrplxESOdBBPT7j
7Nz8BRgQ6qE5eZ2eUkDuCPC3ZvPQSdDkQOooKQefakg2Sv+mUODz5qfaEEaWQ28h
aRv/1sWwqFMDC7aSZ1oSR+tT1/GXosUDnVC/0WY/CDWf/G8BfR/VChrKmqOogw0+
mFKWfk0U1g/F7Pu+DFTJqC8T9zwHJP8WEH9Kb5VtbL4WEOcgFcxy/v938tgdDmoO
59AIGUkLun2vWiZ8q/0P1do8zPX/BQ/+LekdPwC8ppFfVWMqikU4MWwZyv2jlSIZ
2QZLuA+4Zgvgj/mPztkG5wABin+gxMa/Abs+1/A4RrEQEfBdp0Ha96pu/ERiGg82
3fwqbvm5VG8UBDcI3sye+GbVZTvk+aK8sFZyovvW71dptyQPlfm2mGQaPXdR4cAe
bsck/3aco/eMS4EL/M9Jlxv3TrKMo6KHc9Tka773hSl0/kLbku58BYEAZH8GRtep
5dnXzveckVyrZ9p8mShjaXfrip4aGPP6cQovHK/FLXqhtlHmNk1y/ZS/EC/JLmfE
V9tmnfWBuJVe6nVGKcIAf3++vmwQIcnJlCfZQ1Vnuiy3yTb/2jhzg4gIC1vr07ke
voCJuaDolndlY3L60vNzRVdH7OsYKmcQH/eideUFO1tjJQWmqeimZjl1UD+5oiET
IJddRh+4J9nijK5hYrXG2NGe8liE8u42g9PTa2rzZsmZk5wocwwWiESvRnJ8rv+8
kQkJWBQHEBSA5U2wLrG+Jlsas24URaBs7wcD22e/zsP1Z2rVghQQYkUGrqTZSTS4
RIm/aYcLdJa7pn6jv+loymER788VDqHigFp1ZWsAt818yYKuYWU8uZajPDMlgWad
M3cAmwN9ya0Cu+iAL2aDbZ7DwHA9lzN5idOJH2peviuSwlHFH7B0EoSKEhIcVk1h
BkLhq2Prv48ONtPWfTelLpm34boqxOa9Aqafocw3gv2eLYjnD+R/3BRIO2pdukBa
QzZH84kKxmNzwiRaFAr/BQpcUjcNY6tKNuoruoZUymSRxQ6g3Kb/2qu1gYtn2+sc
8s+Jh3CaV3+5L5cGxq6WwEBzIbD8ZOW1j6D5kVtIeQaoHxAmYf7o9+MMJgXiqNAZ
ruT06DNABskNJ+vPGGjMF4ryX1L6DiXDMcZjsjC3O1Pf6QBkEBe7ljeRn5CMiSdc
CWP4cexB/Zd+qJXiz0xmZQnwlQXNtY3WvosM68swNKr3G0UPbOVfrA140mlE1pKk
gDvmJUSqEtbPr7AQo2E56HLUqv+G86bgcl7saXysOImePYvlGvWP5o1t8xhFRDB+
olZg+ZGSPuJi7A7PsmByJgKVN+sg2QZ+pQe+EB9KctNfYJr8W1ZJPc448/L+hV+g
kAmg+lf33YJCMILf93kNgEcFXN6AtTWn99l60vnQIZpVLwfWDYj5Pt3KNJNy/yhJ
t0QCPHm6WpGQI05tuVuO937Jqmzn86EDgkVftkLoasqWAZLkqhimwJuTPZIL7bpm
SieC9ekT2TZhvlYSVCGA+AMTVfWz11jYG37UBom+PKO6bjWWKXn3QizNoEFJYt7/
/AY7djUgywvkcz4MWQEJcNrgr5GQyJVChs6Y8eX1JNHkDZub9Z03+w3JZY3fKm9S
/ix/6iCCvUp1ba2eaXUS1Xv593sv6lr91ZsIcRg1e0Fzt7zTnJW7x53jeGcDRI+n
sYscWit2HfIp1EAPCsei6mRx28gyfJ0nRI2AG59J+dxCsXK0C25f7HJzMGzR49YC
7nnlya+MFd+r1aqhvzKgi2rzOhgvpPn/F7rftPPs/ukJSxcfrrrZIaOaSTEAlDO1
RGlkacBw2QjmPnSbdPc01RRvY7y5a2HZqPV3M8SG1iinF4aCOrilcuolKkFWeDj5
psu6Ux9fCXJxSdNIw+XLtb8/kb++bQtWUfp7LgGfLCBiK4Iy/NxKILNbJA247Cv/
fH5UZxTmFnDNWL9cJcmGI35MvDervAq2zzSYb6ASSpg+MDW+v7E2aiwahIRJC/29
WQLs7nmQ2KAfKjRM2HaVps+rWwmOjiXBA3vf4Qy3XzCsxidkMIrHMQxGuBHhMJeB
zgrKf3eUxEy681B35sXL6HWEsWrzI3j7TNXQNC5TKifD127J79IAZ7PrYHew7AZG
EYsL/WKcQ7Q7x/kPNU230Sh8vigJkhXi2KXs51077Hf3NnfNRyd01dZFqaRGRPw4
CKXwvpNYgth7GDVzW3QzG2o7xUJZJsU3Zf9vqnkilXg4TTpbHSLZ9v9AH7nVhd5q
/jig4PDd6Hxy0p8mdkU1OHOYs5MVrm5eZjwB8RgLjoVhaKUbGJVX0W5IAZzqu9rz
9NT8ADUEW/ufHy2xd9zp/K+HD93ET/WlOSxjHmtTbJIi4D1TDVG8nzpBp538mr1C
wDUobufOPTTilvTFZcou1WX4EK+X+8NKYv7qEdVbFeg2eEUnmdLCCbd/rO2TJjBH
8h7OEbR2gLeru+Y69AbzwubEApf4T528jBxzLuvmonduVHQhpgRGHkUFQ8yVvkGL
ScydBp6aowB+BbEJPewVs96uP6IP9Sr7bCpxgHYm9gt5/nd5aTH2d7ewRa0obd1F
jwhCnL0uh++qj/1QatMq8RRw3SXQBYqLs/m1URLYigi8uYivkhZbrr0ls3ECk9mx
3HZeoJy0bhowdlHDKBUjPbHkZu8I7j05jfHybgYropEQgUtttlUbLNVLxV84yTK+
2C4SGiJ8nBHCu435QK/hupKWiNVTm+sQ4Xg5ir4Mb/8Wp+Vxhz47smsfx/XgJbcW
95DjA62+uq2L9UmS0VZx8AzMl/j7XCh3dbTMftJ0Yf3YhouPz3ZlW3IXbQuZ9zH6
fPZQy/4zSgDLZPd0j6fWmev6D27ohjwjq6oLqa6FfXk9I4tbpFZSo/lMYlO1dHAB
bYkZekL4pi24dylO7sKOFjlyUzNJhY1BOJhlM6TOhZOoVXiDKlZ1bge2h/jjnX4Q
cLO4cWzj9FsOvW4y9+N4Vw+xmLhTdxjDyT/GqMzV1Y4EIoP3fv1vRxHX+rPupcSw
v3N6n/OTi4CXOll439GxuUeFt8Aq6UQ2IjYThwkc83LfAo3Yt4PdmMkXjeaWEGNd
gvWRguQOWvCAb0EcyKZTtrlZ/fh2eeiqPBu0qC2CgjcKLg+/MDxJRCqGJpQSk5S/
9Jgcyz0KZEzs4VKcSB9RU3CRC7p2vg4eLHO9mPVA9c2+5uz8O/mnBhYwvZX62C8z
DheID4fdJvCk67rE16AG6p6flu3QDOsgWKr8CnnmEODqqEdaQ6YhLVIU3O24OaB6
XBrmUCZc13AGSUSGHiLBPDNpeRqUQJy2LWfoTWggA6t2N8ESY+htTt+PnBESedZg
DZ2RGALCy3Abu8gVhgfeq7FNdwD9yqe3E3UMXVVfyCVKHB7ddUwYaMG1H86jtb7n
Y2pyyBdEiURVwZDYrbdt5gQ0FT3qxeJXibG4ndIgcY4mdh0w8ecY3t5fg1VyGicY
P/LG9Qn1V058r46+pxjicb58e+YRZ/b6R7wJURZoN+MYRFiMPsLz05QP5Z+k9T/5
Vkt4JCq+njJ+eyYkBthRfSGEmZuDoK0d4Zk/4FkOmHEWGLlPTOv4caUv/Jqtm9AE
DmGXANz6ggPa/F1RyGa3yBTsu/08vT2tokSroh8WjGdTwPNaBCATfjTdS4o7NOIE
0cTsDjKa20mLU25pR+R9VLGY9h7nCilz0gGhOmzwRSRsGh16AKtAMfQnd9n3ixkz
xbcgtKwyuRpWnYfJj7BJlhpXGlxRKvHNYsXrerCuZRhEBPaC63SCBdOtNYtxkIst
hVOpbqRkr06qzgmRcI5MIO0zem09OgiGtVIWA+m1VP1dHd0qXLyKaa3s0/G6tj5j
aDeIToiUTY/7PyS2enTJq7ia1T+niYlbgsjsNgp8PJrtvl7CZnG3CJQoBMuml3Kq
rjau0BfsyCidf4j0hkxXBMXq2DI01jCvk8I3j4qDDxheBqzuGa/LTErcsmUwRX5u
24mUXLHloBPM4c7WZK+fm3wmeKcFVNCBnfnO8C8M6fyuDW9wj+KAc1X2Z0hCSRQE
CffDNnHC05sYD6Z9S8eyri0xpU44gMij/efbDbALybtVzaGPzJFGhBq4Lg3c3QEs
ZiI5UZpluVt4mm+p8nNelh1VHRuKnFVNGdRmqCut010lEXArM2L5+FWt1+b/VMLN
IjHMVoqyY1wXXKg/WSc07prM9+6zKzV1aa+YAoUl8FZH9EK0/HrrqJZ170QKlO+p
OQLt1BTFGojtseVOZDGpTm9k83qBMF3lvbtl9yQgrnM7FaqzeTcdbNAu+HJrQ+lg
dotTGYvprgJQVwAhdGijieDxdfE/fswchWHSMjOjbPPuIm784h0SIIU0i3m13wcP
ktiFVlgQSGxxGz8uuATdfxFVEjVe/SMX2TpfWsPKzaBy82abQIiYy10JPWDvB3jG
HACqa2zrVQ4nUyGgSzQ1FdkKrnOpgUeLQYGEGbt9xU/wMI/lZ9m71Ye4aRnr9l3L
gOwKlBO5KY0yQ2J6GTyp0SiIEfFgItqBFDCeVPnCR2dNu6X2Jw56q90Ynr4aLzV+
0hMpYelKmEeWyfzA6UuIjr6iw2UTposo7jifsVcul4YlcZOBzv9PD8rADyIf87rM
mZ7zZNMRgxDObpbdBzvSOLojnxp7P4iTAE5CYazPh8/NJpyHShhrslICDy1IbF1N
eDOkhhDwkn2iRtWXtI/FlST5Wo1A+JVCHTC+GbCOGrmJ1uaZAbfCrfCsApIOp2DE
dwPmQet6b9jItKODTPUOwPC9XMg2T1fEkAm/0m1EewupWZPVl40fi9Z5xsDqVqXb
NKXH/cURNq+9qhtDoaB9IcTGw0LOC+bIAJJbIIkH7ucH+lKlHJuV0/QT1OuXPH9d
nh0od8RK5Zo6r5G+HjBvX87vYl8lNCpYJXAJT/jEvfmiiAJ7CY9YII81bZ/jJ1lV
uW9fXA929gt33AEllWRfodN9jlJVTnr0et1KFtvlF97ermR1LYQCZenOOQ2R3nkg
LieYyE/TFUio6LrLqIY6lILvP9c3aqGhhpbeSNAeo91sMjx6k/PV/H9DVkDjmWKf
Qzgfk8+LOvUB/mVJmAnPIBF8dyBHJ/qsPB1uphSTYM2JCGjyrjluRhvMGG21wSUP
DSAU8P9IwB5IJW+LYOBkLPsRYf3klyVV4ttmwXRB9rYnKv9PRIJKY3ftW8C9UWzZ
duSUxG5IuXWsF4DeO7uAbjVrZI2fdQ9CNdLFov411U/BweoIJe8WJ7cUJVNC88O3
wDxk/Mv2eASpLFwVktDquBNIrieYFCLURT2EajvlBM8TWX2OuQwHjtCiKLZYEjBJ
h0kaRW+Orw7JoE90DWJCQCtxttf8RJX5T/O+ju6rwbEal1bPjoswsJNKG52gZsqk
+yO6K7BklfYZiwnrErMckC6aof4f1GB4ZNfgD+9ubRqpkO4dp16gmg/i9cI6fxeQ
8wl3W2XBsdOwawoPOUkb5jeSy2uO3mbeJzwyYB4kVzsOJ8VNXJ92X9nGFjVKZItF
DmWmApIlx4MiCexsAeDz/T8gqo3cPzm4TUc+V0S3+HHK/qtwfF9QQzWjXCARMH2w
u+RI6geFC+0pTcU73jpupJS4Uuw/GIg6vKRwwAWFSxPVHwjmjeaRKzlnP5jds6EE
0w8oHcStFx6LUN0jZCYuVl5bx85/q0sLe7b40h6SpDur5y3hb0dV7BU9dciOItpI
0XojrBerVWDnjCgT/egeaCucTR5tk4NyDcJT0cOlv2dhqyVgCaBdVbk85ap2rlJi
9Hci9gooJA2gnZVDup/8zrLobPwAogv6oHHNs40Pr1z8GbE6XZSPZaiObjTUMaRF
bBqgLRTkCDID1F2cvhfzQVrf8Qhw4A0+KpouDQibm+JNKmtf1PBUVTYRCfUtEOxR
1iOGaDQiO52vwvI8+LVnO1A5r/D9kXQrOfW1bvRGX8O7rvIg2qMaKzfQpfgLRqwP
m4EI/MtjahjJw8RChzk8KlbydFsEQ09hVQ5En0r6otLm3iM9SFxEvbrCtic//7Uv
1eeJMQgnRqnxEcKVDU/pT3kgT9CoV92akEuXiQJ/KISsUtrnkM0/ScvEOUqnn0w3
+MYbZeBIoiLaHQSWrt+0xUWMvYxM0Uc8KVwii/fgZ8CQhKzT49kxvSfq0cLU3/Py
yF588UnaoRpLHFCC+i3tKytzGSGe8uCLtOgbMjeV28++zbCQMKUZtTdqg8yAwZzZ
2Qz802WIPfj8xZmTl1Whg2xS3Pqh54GZwkDAcyXbZGr+uQy7OaLTqFIDi/JNAMUs
QgudvXogOrx3N+IrnXfb6/dFAjCYIHq9VLEWMz+TAH0dCezxMOpip0KDbZiRuIUn
rMAXd1Sambhx7AK/HO0Ma3syN1G4OFhuaucgbh9QDjRFcH8/6vxKgDz8WCZ+15cz
5TXB7Z4lPZ08owzAmp6ub3awBXg/GOWvnAJuYYGu9thqZiJJqjzkL/qRm1tQu7JJ
/xpgGIK6lehhigxAMaG7frCEjjQ9HPTZYOYgWLMj9lhDsSHSBSueGBSsQfB+bQFy
n/fIP4g+frfB6ScbChGDsTCxKCmVgEUTL+41e2bRO4RIIfoC8PPw338jZb1tRSDl
x1T529GQwV3WW2WKC7hkhvRovL0x/BOuQ+6Tox1/HfCUI13A8O63Ee6YCSPR2ED/
bmcJ2YkZQCsQIbLFyNQWx6F8jSUQeh0Q20APjyrmvRac3Y1wMt92+JwY2j3nTmvA
BhMYYfLGgKZ1zB0/hBXi1m+Qb49oTY66q8KQFaP0m7i6vyY2oUDqimwWyCYakEXo
w6n30lGstQstemORR8LwhKV21AjWvBjkmAGgs+Or7gCpe50JGTENbjf0hba+ICif
9Y9c+4bDcw8dSOEMQp73Xsz8ehs2edKFHIWBLzwGcH4ZsucHB7sjtn422wZTCyZ9
TsGDo+xqCXwCRd2tcyU3SYJo2paCoBD5yCQ/9KoKdxFZJ5TMsp6lhi/zeLXCcovV
mD2BQPXIq/UflKDM4oTqUhYea89P+X+g25dNevl5Rp4pBtsCgfjym3yLwSSMs3u0
w3h3JJD725TZnWhopIIb7UWe4wH+AoQZ3OtfU53JDGMff/AZAJITFbivfG2OnwAR
P4AnXIFCi957nb2MKMbqmLg0i/USplT4XqJemug4TSS84/e7DQSPpxV9ucc6L10U
Vhv4avbP+FTW0LMcVpcoy36RiCGyUKpBzITzVpQtH+7loVGJ7PcrisdODjQmEDpm
HpuRU/IY2POcecVJ1ILyNalNjagRb0IcNhRnL/sAtknIgi2fmzuEI7xI6fLAnu/T
Iu0eziyXbfiSb4q43MN0+0aRimd3HEGbkZXPoSacmnEaoQRlM/5oNaxI1AX54xJH
VTv2q71oQN1KE0dxSB+ryLvA2c7AW0bV1+LdA3bDNkuwuevFYbpzvr5YBZtjmsHB
G4AiZbWz63tDnHNzUseXn1mLvrmn8Ve3cnqio8z0yhPGM+2etddBN8F9EC/Nj35O
p3FMzmt+lv0JJXYm0reI5hK1Oyu8jg3sNS8uDCfiB77dZWqEnUTNeRGe/wgJmINk
XXN4lwKfXgyoJdodSTIYRjwHZI99Gy7ziPMpCwR90fOdLXupK0xQptPAUIvJAH0Q
ZoXxMydNhcrkWrQLIbL3p6JiLa+b7npIBg7EZc8C4Hcl1obAVeiasD487gQ6r3Xo
fHMP3elFdjZxZ7zqcsaxm9FXhR3yhLsLyRjuyszs84ekhKVeb0JiIMcW/WkuFm9Z
MD1Q1Wqa3K7U6cyAfEbqG3HBca5OvceEPcQ3Xbuw7F+n/K2QBiBarc1Wp2/n/lP9
1LNKUDlHSvCBa3IB2QsC0yn/JBbrQ1U/sIYUY22NNyCntRist8IjAE3cboRI5HGS
+g10mAMhvvhdwfyIgjXbLQ+aPsuER9/0PNzUf8BqUfVMRSxNb7FsUg2rdVDBHxYr
Zddry1/qtZ+WEcUDXf25RR9hqHiiib3OikRN4cKbTcJs7qbxuR1n1O6C953mihoO
Ur+RdSCmkQdGszwW3HKbCTuHpUq0FOD6IIoroRzS9YtbkGeQJ5A9xrtoFnpYTPQx
MuU47/tieiszMRcZsybNfjT6+p2ppKpV+utz/kEYX0TgfPl2OJKyfyC7xW9MfFUQ
01g0en3xsf+ujVweuL2WbiJIBh27sr3FUjOka9+SyOI5c3z/0HkPSNe5/+kfYWKv
AaG/u8Kvpg3EvdRywvEhMTjAeTSMy+0pHlL9KCAEOhlPZ4yKYyHEiybJfxk+zumD
/oCRckyaKOz+wSwJDpR0TdTkB7KsHCzHo/sSc4KDCorZLE7uBxXy2r+P9wWNdmuH
g5TqwKke6rGmUcT//slGK1m3gn7XSdZAQDICoQzu9YiSc1U3BEI5M++JnO5wGA+S
heB3T6rViPiGzGlPTz+R1O+M1tsQ8qUyDM44T0E4AxlYAVyCOL2hy1T8qDhBhqnq
0TQ4QpL9+3OKJstSfGzGmmjjkdJ66YQ0s6UurkWFS4ZSlFQkcf7IJhl/pAKoGfMA
N3Wn8yTAunXPPyV+/7XhitjePGVf4WoSTdSeMl0U87TfMW4PQbOh4Bon2AdD+XLN
lg677UQSjJS5bpVyR1Lfc9phnTx2DxYlnyjXUSLVIL8862hAsGSGsl9ie0A+PvM3
5lxRZV+SfKCWnRIp2GrsnqzXmGXtfKK72RsapKZL1OK0Cvy3XBjH64ikJ0n+W1kc
I1CLLYzEBtIHjqBAhWnkGP90bGft47VxLdAfykK66eoyWHtCNzkhwHAHyTQoBhCO
DrMAqwOACWN71A11PcXo3VJ9guLBZvFcE7jsaIXn1nv89uK7ziDC1MoyozfxIBj1
CS6KNT3kCzHMGyYn4J5xZtsgBw+0NKPUmz4bEvgBTyovmVCppL9a6GksP6Rl2pU9
dPxVHKtAV+B12Wfj2ECTK86LNxrxEVXo6c1HLWjQ717aKfgohHAPZgse5B6YKaaA
OTuujkUQV+Tt0ui9+zbC5FHNVzoSYiERPdBPAGgWQyl11/jwppPFDtLMwTdS5Qr9
1JrsNpGrA3Sy8lmi2nenrR1xJKjESZ4uTrGWPyOmsU7VfR14gTYkRIU+CnzatmMm
lx2Pf0Sbn29XOlEsEqMk2jsjFx8ceseqyXsuQ5suLmd8ISnL6L+++qhY7tAv6YG3
5ZkH5NEOEQg18bv+RnNNGwtWi4oABCfAqmrMBL0ItfDO4tzQpat7+BiSGM9gozWE
0WUJdAF17meCgdlEH0WAU5u3tlAoL/rTZfbNvMLKbytoFXDgjQpBIkfxpI6Q98FO
h8+SNdGDsGFBw/1hXftQnJVyCTGtTeCh0/k0HstWZTSfs4k2ieRubnOShqDhFuaR
gKfokp8OExhumDqn9UwJchAyHcFPE9MubpsM3V5ufscZXrWaHJVv8N4IQ+CNRsPL
dapR+RLBddcqI4VGM2akBgHhYxl+8LtP1Xss5Gy5lwrpyK0ir8hZZ/fOdYpkdqca
+hLH+rlDJY7QCEsw6kkWHRCMlzyT3SkCJcYMGgXcOdJnmEdyILCJdJjC7CNslzm2
GHYLkDXs6/dm4qV/0Dy6ykjQlr8wwQB2Tv7agDnkYRualx5U/vbkca+srG3pfz4D
oN7pMG2T7y8McxrZ8LW8ZZanXgPzGrjKhQWEXY2mnCJI4pjeAS7TrD5oItPwUEgB
rqR7iu65VGQz3rfdJsiV94vij9cq8WRhEDQi9o9rCT31t6ZSfMgbR/XVzBWVozrL
GauOMJxKtVhtwA6kCWdErtL8ts3ICYFhed0al4RpS0OUFo0RNZvPktsypbd4/fnU
YSJ2vcTsgawKbKu7TX3PVFRGDeqNb37e2JkaISQa9mVMQ8pHGXjnTcoUrFPQSf2z
qi+8i0SCfTzCepEmc3BbEW0yhFL+Ml6mZobyFYwsiNfdgYJhoNi5HYIVwVtYk7dw
wx1jkPwjl2OKUybBZKNUibEGym0RftdnN/hUuS33UZ9FzjAXl6bHpqB+IqZd1GVa
LIiwytSXF5j6kOIjN2m3HJlPZNpQ9Y3oIeIsnGB1LIrk2LFkCBWiZhr+1iUGN5fu
7jJysLuCFtBPJ4DvArHoZP4npQFCUx9RCQWXUG7p2ZTWv/fr6TSg8xBNh/qNOPrI
IBEp3BtmP0vkCqoTIhXl8XLIHP688vmjmhrOZuCUhyOxsYH37LUEBwupc8Nqodpp
pculFCn68IKtuCkLSNsXDaWw3AyBk4lzgMxcF4ePAc03tFJvZ9Y+ZXLk05vsDgwT
xOkJM/3i79BmWc+8YkCmc3pVXH7CnOILjWhIdQP3os9myEJKAkN8lRgnCv/lsJEy
jZrIMxDSl95KR+9pm4WrpEZY9SRHGR01IZhLABFkq2mC6/HZNxD6rkeOi34VnKbd
ql5eEnvQipJ4AyTzCb9fhwcCmd7lwo1rI/OUxRt5HFVqHLwoydUHSU+m8oyrpTkX
CPCkd0OIB07owYxwzqhY4rZRnhmzHf8aHz7dXYQACHAI6+AqjP8yqxnvTJFmZ5WZ
0JUtp+TpHdavwzli+6B8hTNPkg1ednnk3P8zDDSp0kM3P3H+x7u709dZ3kt0doYE
FYkpyts6GdN3seuW0zMttV+7PzPOtceqCwJ2nHzDOXMyZ0v6bG3wHGbYepS1JHeo
MZwAgSzceVGMnq37BpJgPaJ43WTuStUlTVU6sLpk8y+XlzyoG7nhBzsqetQpqdy4
0Phx0PhEMBu9ON9bi7+g1/yZlUj7j/3y9l0k8H9pieG4ConqJfufM8KFC7EyvqnV
oYc20LT63J/jFsBRwNR27tH2Z9r9/+Xtu6NrBaM7Qi9kLTe1BcuvPRTWupkRXlKv
sez6d4euZVWD2KUIJXoiNprg0XHzPfCzl4VNk+6/txIrARS5gDFS8EUD5wAhOBRH
jiqdhvDmZre/VnIA9pNSOlBy1LVfMh9bCL+CT/wMUb4qfCWonRqBVovgWAVIKJ0k
lJwQZRY7K0iGF/ejbISGwoL92xa6ZG2k5pD90GRGeZEJicRbaaob5dtFvuZARMnC
y/0OV5r2H5Q6hw/faW+e3BjKZxZUBXEcTOrmwlsDe4zVrZcWCSdlmLdtFTOsiMKs
dDYnhlxxykB1pZTSuNJj8sCJiMgDY5NbQILe0DpD6/tfQI0OAJZ10F8xV9jp318k
5cVhx9W07BpP8u16iX1hfJtjF3C6o7FXSBDaVcFVNt7s4xANsfIYttRq4MM0Y28l
WzWmwYdJFMGUGQJgbvTyCy2AyTVEky1jUtTh+K+B3xgK2zT0D0uhRnBBOtgymiiO
y9GhalTrtYxo9XiH9MhCsoiIEDRBOkHraWCglxKIWUXlWKXMQKgYd6jyqp+AbWSy
bvGreHzzf0e0x9RNA3Vl51wBQCthj8uLWt2ott26QYcrKm9xTc6s9411ZlZbCBJU
sZRSMe8RreqqOv59PyBKG7AalW5JEbeNRc83yNHu5Fr2d5loZR9gft3TWPI/4jfV
CBjGYHj2hFOdGVdatsEzb7OQXXmR5mXNLrJGbFDlr3EW+GQNLJFvf1CwSVyVRLDr
V476zgO0joE7oC6cwndEz2S0Xf3HDhxakmCm2UhbsXR4VYNZUcxp5+uokB8S+Oll
F62mIYx6KF10OMoen92S0a/MBknFwbBXR/Q11wNF7GmLPe3kVxrV7E8EIcWjStS/
tt71FI2yzFI3+wFp346YEob64lrNH6/g23f/Pi2dunKzLefC6Lnbry0yeNewY/hN
O/qmZA5z+2W+0x9G4V3caOQkKRd8BgJcaeYIX4aYwijFa/ZJXT8kuLCuy59bSUPd
FUc7jL05FpKuH07bOAMhZD0yJSfeSSq/JCZgYarMNL6NjLNDMF3X/wsJj3/3Ar4Z
TZm5BWrJwjmv0GY00aRcGrSGpSogLrbjwA0agx+nXDrYzJbyI8Z75SC3dpsfdbV+
gc+NL0E5rXskzPbAxsdrYFRkeWq6TeYMs6zn4oUDHla5TqWPYHrPDplIouH+rKFt
1kNUrxbUpD9PVUYy0Cuc4sqZavuI2LWphjRokLbrORwR9KM9sJJ0ChKhhUZgwhzM
fMJx41bRumkHjv8aLZQ1qtOeO2qIj5nJP6YZV1CiO+vgtSieS/wHwgrdClOAKN3Q
98qi52pPgUfmEuKviyvexcuJZ63EQACwOD6EHDEx14CeVxM8wRkGUgE594xYFh4e
qaqz4upwVexyUW1iCL7uOufG1BAWKiSXt47JdEhTAeEPhU+UJzc6/9JeNd7Lgq1n
Ob30c9MeYqM6fHaMoeLU58yKSguaCa4YYr4ad/NHWAe4ZBQbSX9+3F8L7BreTPAU
RDgz/Jy8fl5Rf26158mkK/V3oijldtvcViHIxcnElFG44mwyTI8CWHCYUJB2mXOw
wujuKTFx7RyEWt3CcpYJSO5sTExIrZVKaH2nfBmbcNKKeIYFhMCqXWIwa+YC7Eim
VqSntqwJULO/MFKXUpY2EE+ZkfDX+gHZM3VTTsCU4XMqweIeOpod8Z72qb19r6zb
NXeW5ul+yWqAjA8ga9GCEmYbOaxEzdNTclsXqMDMGnLErpsiIivbsm1bh+eg9JWC
s7Lds6X95JISlHfRuleiiy592sTTusbgAFv4J3arJViesTf0PwaS4XdiclpKwXlz
TvGbiSNlRDl2UeoQPgX0/fVNCmkKDBWFEHw8MZkBXHpRUl9QVrtuCeRLQRFIjXIa
wF2NpWw4vFu0hFnJobsT/XN+qrEJI5k1WCQ10zEug8yWyj6NWQzwYQRw1C9OS059
5tLo986kdxm4/88JjqPUAN72DFQp7+/hMgWj/HRm68dg+XYFqnuk+jqtdNSoBtVH
W/ch9+ZDIp1BV21MqU8nRtF4vlJPn0grREYmHH0TcwSr5hr4UjPm68LpwKngD/Ts
nVsnmVvRN/emn2iUS5qU/e8ORgZJUYDL0yikZ/gMi0G+B7oqin7qSLblFKm8fF6m
Y/9Yw4/kUrxm7L6SMgTEK8wry4XRo+gpFaYk+OuRgAlIy8oHxJs8JSprYJiZICl+
TFW9rohlOozGFD/M+79JrmtpJXfEuJJlnha8ZwqJOLpzBB47ScQo3TOwcl0WUZaw
f2N+WWvyduOkg9cFdkkfdzgv/0EFOQNpo48X6d3rkwlizvy8op9I2BSu4aX+6Yuq
GyC4nxIfDxzRs66EldOmW3FnTqwp+r9l+3bv3UJHRUjTt+xgc+JiIJIoIBMG4ACR
x4ZyOaWwvd7t3ZRt90A66UswVM035ZAxTmnG3PA2CwAcq1yc/FQhv7UUMn6wdCe/
Bf7v/tHQSvd21hoW1mmre2vX2+dA4qS570/Iq3o7NtdxoLyQybTB7qxxigqFgoA2
dxPpmA7UsJZcNzaVoOrnSVFMpqWMMWFBsi0S8PNPZXoKjjRJfH8FWAE4sgNKFwKQ
j4+F847dGJJnVc6qmpRFg9Qy1Vr6mv7sgOVSnwhT76DHwEI2VpoKzJZt2vge0qYV
oI2DnWbQr/qElJWMz682yG0YveM+eJCjKVyT/D6FGjsC1YjBmAv4QxZbiWE2OQ8v
JgW3xkMTpkkXhGI2HXvOp7R7fcwPaHSUtrYCFMiwoSfWE7R7smkF6f8pUO6oT/sL
k9CTnCxAv2pohanATq0vrNruLYdSjogingCg3frpVD7E+26ptP1PrGIOrKQ+lY3o
jppNJ6+RB2goPPNDB/gqRlItgYqFAa2gQZtFilGPnMLTZ8gKI3gYlLTOBuZlMsJX
oTEst7Yf7r4QmmMua1BCDG1z5SY9n/hY/3Ze9JLiNN1/n61arR/ZcgKGgNDyWU/K
qPLU/a0AJuLq1Yn5XQGFpW61ic8hIhbkfmuf3wQdjwpBPK2fcTRotUi6LElF9Bmi
MtR0e19rorFLOd4RmAr2fvpI5djQ+SQyX9A9/QlM4pg1nzXEcHk7gCMOx0vOHsdL
KWvLabK/8pS4kqappTLGUrkbuhV8LZ6yQFDX8Tnfoct8agkLqDYuaVabanBkSsoK
E/mXbw4cN8Wd51IahM+vSwf+EGggFKQ4ipqZuMdDKAGeitNiZ8w6SLawOTHVA337
kjAlIizW+1Gh9j/+NJZImuT0nMreu6WML6QVEaxtI4aumaC5jAVu+71CTe77AOu1
mWQbvhspouB2mUxCePLULt/44WP/fEpDhKzYtjZw6bZ2YHvRaVvsaq/uy7lu5ajh
7xF5ryjOShgUcfJhf7fJbFOezcSq97fAeho0MLf6w7VCodQqkDUqxy5GBny3gL3X
dskdEQRJxyFeOTGBEbNoa2/HMHmh8YS1PdYGDmo7ENbr7pKN1VkrGSc4n3wyLSu5
aha8TfOZlgJ3MbZBWxD09CaupneBI5BAYtXlByCcgs9ooff/g6fHgDRycKpBZQ36
j68QK2To1rqwJUAT0x+U36H0qX1DCUo9pNrhko3A2kLsG9EmPcgT19mMHvgmDC/u
qc38r6XMgBpLELi6URvuIN2eDa7e9GxAp7d6hnWSd2VBV174oB8EA6fPVsz7Fswf
yL7pagECmhvfzQxZzMqJxZ0AEHbmcANGyUY7niHR4tIh0zTRSWJj50EcrcmIE7Le
BftuZXf8S56oV/+W9A6gdM5zUOzXk1oy8znHZz9jzcj2Hp9UszN1bS3A1BQBrzyV
FYdb9CaMw1Lu65p4EqO4TnfO/fMSREQ8WMqpgs78eyXaGUBWsNTNzhDS7C+38m9S
w8Wu2b2c+Uzzvw+2Ic4q/bGxb4PpMDIzeZYAgJIOICozj+7YKQDE2l52uQZhpfVj
o7ja7zH53y9QkH+MKog5d5jIt5okRRZ7A1kbdt7bpZOHqhg2M95U+zbgOhRsY7eQ
9kPg6vfFiqSZYWv6FkBgBxP1QhBrDQz3p+nXsdUK9XmXXtM8JzUX4EpZiXi+gmTT
iVe6F/Q+ZLDnvERNiDUK9zLm+gm2sHFLd9aZfXNr+5zVEjv64MFGf59uGUeIN1rr
RT2qH5hZx68mRaNFdJGAFZRBJWWiNlcBO+20X+gWyszBwb3exbkXKnwXVvWq3u0J
ZIVNcLnJIFieYiH4xL7vhPjlu8ZkGawokiEMamldbx/pEKRshyi+iHrJdkSP5n+J
fwkl8fVYxDH7QuEPmv2kyaNFl92sWr5DqG+DwahsIczm+9B1hFQeuyIVbol0xlGO
64/cbEyJCeVB6FcqxkUUhpGPwFmPblLie1cRh03WAWD3oZswiJS4Dkm3yXRzOXLK
jVYj+rFcPEqu9Bn8OZnFWheEJLjPZy+nQLH+ov6TZMwyxbH5CTRrlZ9BD5PUrlbT
sqjJA97YnUXszkR33P9o/WawKA5DgVULrmuwZ5JO8dqld6zJ1B9AFA1ghiSR078K
lIBnziPNdaO9mgVMpl4GEoOHfFelVfargBOtHaoSzH8csouaiP/mH20HtYWjuEsq
+5vXwxeXxZuG8jMcSyRzZuO3BZAiji3DL8BOShUszwS61QnkaReNP2UQhKaPJWZh
G0thelrHIbyj/BVycbdQqyzfpZL4wx/P6JdGONgf9QRzXm6aSf66cd4XI1uoAR9w
QoICIKNhzeGaVwQPM1zIFLlvKv3g5YHS9ZKfjjMPUvW/dfa9UciwbnDD+Hac3Doa
imO819HfTFENtTnrvRoMymUAwWWsrBqh/QsEymztWBUAKfPqqvsSNeTTyeOvAu8A
lTaVcyxJbnvzLeQP+5m1RZQXJQb4kvMgh7PFwpk/p4Q5Cr7yAakGhjnjWbJZlAdu
bj8VF2VJoxeR0XnXOU9wTKJKVfqj3JYIZljxSth9TNBx3+a/h18WIXHutPXst1vo
1DZ3g+09/oIlMpGk8y2cuPC0dnoZR/m1Pl8X86uCXNhrwvl7clmXcQXNsutzQnNg
jU/Bl0OsSEMTinh6v/zn0hmdvYknLsMrTLipVTqc+w20jpt0qXgZW9mDyfW9q+Ng
GosOMu6ZPFM/enSAnyVkSDxMINMmFMe3jYm+JGfQRG+B1PK53xFEeeXg6KS3ZdHe
okFc45p95MO6RKr4Vxp0HRfeXgvs8sGku9reeCZW2g6M9eNHCuwUEejMyb1J0CxG
rLrjOwV9VXd5e9rUB7XUEmPLcqrg4kSUQMaD923d4px2gJUCNgYyti7u6nxbLhrQ
n8gmGm2jnfzb7awKG30Ehk+gphfKu3Hwmx7KErpgDb+zWfXyfiY0i0uYHp4rHmiC
gpIo680KlqgLqf7EMYiVoD8tpWQ00tTbWebv74bqHsUBTShFKxgx3T1JMcqg2ALG
0jOk1pNCuX5gmYUNg6WDowRY/z8WoDbHO0zhjUWIGwwCDqYhrSFTZVEbXeGtLqD4
I5EuNmN2OonULVQ07xKRZ/jUApW4vNnV2DVq8gESHq29wzHwYuSuIfrfeKTNoBYQ
8uGLjvyFeLBgnrJK6+z+fFVSop3FvKZvTFgpOzMfZtfcwVfkO3rYys1SKRY5cLSy
o6FZeDrV3ZtCdpTABHbYfQTxua4tUViB3ocnmiShBlSNkN6gdUh6s4sXrukTbKms
uhYC05fzUvXF76TW+fVupFJCxogZhMcpjB15iUGvxzYOIja4mzMa0pGfhYb6So9b
ud4DSeDRR/Ta3iKUW+oOQFeQolBDRjGWgNamaNcuTwEZA+HJ4IEVS72NhKGqIgj4
OlDZtanQhknIRDfsZZsYWdmrVp7ihBi/5ukWE3s8iXmUEtreDNp2hLkwCAtL1xRO
Ue1AWEdaR8moxUePM7x6qmuheGCeqhrcgRHLCWIIqQxZ1bYYqFynkEyGuU7gyXCX
ZKcQ+P45/j8ksgf2WRt6AlH6vLGOPqWYmBzUv8Vi1kZk12yNxE2ZbJnRZ78QP0Fi
qXmXtUXocFqfI8vJkiZa6K7ZRrKjImj/G2EHC1boZfsEDgVQeljIoO5hvplLiMIK
C3Q8jNUvn0eMSloCoVpnKULAy7jTvajVqv4pU0gGStn43f2OWXbCEmY0Rnv+wibO
hOwszSqpavVWP+ER14ZrfuibqUgLrk2c8PbUZhMtOa5fOyW0gwHJDzk/6JMSDdX3
aa7h6LOWgjaxv1H97YhEIXM9P6+FbTv7wViNKbhtv4N/nUMIpEEmP8n6V1euCNvb
+A0T3K6V1SsMxlEjEISvzOsNqfeaUFc51idfSVzKG0fgiiiC/jDyxTB8BJ7u7pwl
Bh5DkQ+sRGomkCIl8QPI1VaWw48BLFDzMaGsxaqcP8NfYS7pPhiecDpGXcGa2KKo
+Me+NyV0nkPiZPOhD6ZJyred7mJzvCpbTUt4rg1T2oVVjZCvpMFxc8QeKAtQndjI
DzNB0qrzQ7Bnl6Dlbqub/jdl0yeV9/odo6ZGxj7ygXRn2AjcsetoF8QNa2GeXNLT
2kZgRLdDSp/WwN7y/QUKp8NaTh0PWU9jQkkOPqRyGolDj9O6NCwaPli/nKxE/RBx
y1uBoG8OdxYug9CpjyBlRugWi7Om0F3J31PEhr8I4RRJCBmEyEpm6GioKJLsC8wp
pYjZJoX7zrXcwHthfqMglWxGAgzfuvv1YuUK954LgaEh+TbGCv8yC/SZx6eAc5uz
QftSVtG1PMPfZ05OrtdwSw6lnK/u10ITOWDRfYpbYNuy0Jr2r7UQJmlR+cIcClx6
s5WFD2d84p3I/jPGi7ZXmq555t+3bPIYZzviuWR4Ny03D0oAtjSZOXyhCgYIJ1qY
Ncmp/FMl/xx+oUguP2mtxocAxLEUX/Rx5k3PQfmIwZuZO/UC3FCI0GR+XOpyHHNz
JK3bNYeZVna+QwEt1Vru/Lxo5quvtXmrfFgaCk56o3aMMM3UVw7j8KlzIP1UEHbs
GiwvW6CPVRDpkernHWNiOxWSRO2SgewMXaxrTAzGvG+YSzp5CHGDmgxsPgooOh+V
SvgLuQwdKPQ8vPF0qEIBv/TiUJk4Tpzg2JY/8V3EcRY1YDqncKZALcaD9W9BSJWD
SuAct85D5DoPn2do1T/fECGLfQkl4pv6ebbQjxjWCQywIqM4tUW1qMoq/uOjBqFW
RRw5XDzYwb+fp8C1Go782MGXBr/QjbPKa8aiPgLr3iUBeDUpYaqr5UiBfXslw57y
oS3YPa2oz6AHFkUQBw9ApstkLXuT8ggG9haVe/KUaDQrSUkbT1Y43/5uv50F7sO3
1qo/ExRiuwOIx7j19ZoOSIenGdGyrdnuAF2kmL76Zb/EPQIqBs6LCG4/t2+0U9r7
LurOEMyVRvMJDldJ2+ZfZBJEav3vIqTYPH9PUURSZtvaZACoAiDt0ne1AzoT1yAy
TmZIEPM5Uvrvz8hAgCw661/Ht8R8JMgOCcMVIKTl+6HJtzrn8IlhlKf+cMz9XtiF
jPpcve7Oaf1j8fsVIDGfCJPnSlamPCQZ4H5Zzn47rMHduqoyzhlOsmgjbxqXPywt
BBbz/qSIMcoH2go7eHQHkSZf+L1WeRzhRFeel8vW4WIlcR5hZdAyhlHVLw9WZKO/
UT28boRoRDlM0n3vBPdNPpSIUsByZIWYo9EVLDIzFtie5m3/idGOmHwKa2S/xZFX
oszaITEsv0sJ/z3A/Yhscw0sCcbyXUEYC78FvjSPV/BTDURXJH5iEgcIrcXKD1Fv
0naWmR91DZWz//ZFeIiCj8GekNIkm9T7FuldIxBnhdDwGVRzC/EZ0BjtQvWb6da+
hmhBkNKovFm4CSRYMy1waNKdz56nuBNwFl1oSTr8NdT47hB7Ph5TcD3OB6EasmpD
Afu1xDHoN3rydel3QkOsaWid/sDOZoiaElnEj2dmg/b7XToZyxye7tgK4ns1o+zP
1HcFjCc+81gniTX+SdTX6O++rhV3Jh/YrZtw2ByIo9844Z+S0TUwSy2NjhE/zO6+
tV0iKOwhzHOJZeZLCusufJV0eWsLZ1QK+kXg7PamYPQ11iIxB90zqZ+9FJdQTsp3
GpyKZTgdWu/tYT7C3LmYthd9SdGGbyL3HeeRSI4IpA/2UBpHlG2mPakPCkTKtXLC
Bfj9vdtaaTadsfNxge2B5wwv+DJQAJg3+V2dHFt10Axw5AB4op0q91kDGAi9pcpC
PK57ENoNot5EXu+Vcp72ItbGWMXbZFj9tRtfTNTry5t5mZnNHE8sFWjeHA4NhQhR
lFBo9dCoHRMRumFsUaELJEjOvWYc53IyZV8X1G3XiUNIsaOYd8NGACza9KcLrbuA
TVnS9DxGIe4Vtha4qNsL3YI3NbBMpUhKzwPo23YERPhudoEE6H1AoPaPeE5Ova7G
7QFu7LHh/IdQoxR4eMwT7/SDPXggv1FIvu9mokX+NaE9+gdIc/CfSOFEPw7sUWeY
a5T9M+GskLUwHt+pPpCH2LZ04OqSb6BwuzvUW9+wPp+/A7GbuDZd68CIn8oybAUw
VJSI1XEcA1EfI5Bx8ByldDWY0qDYRdpmyL/mLj7DdRScA+IrylZMq2V59ytVDjRt
U6sn4DmGIsA4iU26m3gXwFB4IfixGGBC2olOcWhMUDDjcvPEb+iYhzjRAa4VCmPq
PUkLwwmCMczd0WklO3oIEvN4MFP1wLtZG7kX6ZIaDPD1E/An59o/tZHoJN252nce
CLWNaDJ0fNgTOAfRq88RedmTti+f6NrzzgIKbL6v7C7HdBR3F+oong6aWrgFhmrF
v+Ac0sJS5tG96w6+LkxRwkVxPnFs6YGsaVtFW2vnWOu3CUkUmR2btBy+BcNXiGcr
x/vWnsoz5B6E431YUgZU9GC1mIFwQiEyiZ7doSaFXV/DA/UNrcQSOaOxr5KLNOV4
ZmCx5r4fHxUK9zjsQsSuT7h8SLmt/+YkZmhEF9CFVutLgsfpDk8a8KD2lIxIgbdR
auJQs1s/hlJTVg0GumvFP9qphVF5Jd0THWz1zpfAIlE0GQcGeBsWuYO3RzR+WU3J
zAvOUZYomDXQSsY55pJJOJxOxv05eY3KS9gHkpP15BAoGyJRKmHAeyTV48A9ZyIU
rEk/8ataraZgOYe6v7jRIkYDD91kf8Jl0HM5JpPCQ+6UApoDqcHd5JSXMyzo6TuZ
G2r/0E70aYQeRXQ8CTYEFw9yOa37TL3LEnadY9UYCZzIqU4dC1r+pctiMX3a4lTA
r7eWyFXGjMupzzHSjtxhy+k0bhtW9qbAp2bAOEIXjrlwFtJf+kRPY75Dq5IY3G0r
KWfKFOosf2ooqtgPXVbJOnZifvTAyKDijX7szkQTSBbVR9gMDO7sXjHd4n/+Xsq8
MVWSmkH/YlMPz4O0o69Qdzr8CbRMYasWw1kMBk0Wjx2OGzFn9zEkgYX4pMdw9SXd
6WKQ2yj0v7rofsegwyfqVXIliVWjnNEht330TtbcCA5nXaK654Btw4KbkqZAFBik
IRYzIBVU/gGPRKJb2HzJP/XWiSsDoLraCaPdxH3XmfrJXxdOkWY/u1/1dsadjl/q
jv0vdoTRmeTngHWSlhkirNE3ZX0ttUfXhaHpPTXbNtDoQI8HUK7gmrpwNiQgfPm3
4GU7GKybZo6Tf0aA6ELqGhytQA5c7RPlwjwPJfJKi0WWk3dlJEonr43gLPGxZRpF
cYYBET/P83QQBgELeIbORCf3Z1GOmkTaxgaselk9MwJV0qpQDfD/Y6T0s0uOpb16
FfsHoJornLsTmv33DPindG7qxb0hx7HpJCXmw3f4Q1m2USrITqD2B86ZA3O7p4Ui
tRnS6snVnumH1XZOVG7cmDaaIOJwBDhpEuVno6f/4r9NqJmdr1UikZbZV/WVBxr2
XTMImNPDlpZzvgfAQYRPYIKoGLSRxlElSRbKkJg297Gn9Ak1iNArHHN9gtl+3VUp
ZKADJHrA2CJ5AMj4nGvm2oy0fWSIRsK2kAZjrQfScXSRmj0ZZZD3v5KQpRkIKsUF
nY4RKy7OCe761eVuTy+kCMRwC1qFNf1DtLO9XpqCaIFEsGP8HygllFF8MWVRlHsP
iE2KtNPt2r739dBo8aU9STE8tb3JvT28bxW/LNsXBINh+h9NC9Ncwvm1Zg43SueT
58ezCUdF5IYJKlzxiF2Kperja/U2zzgDDkKafOizph9rowA37SOuSPON9fMqM8yF
EFLLC7D+HS7cK6dyWFpBfdGztE3pOwSN7pEII0gJ0WHixKhMnvitxDrLSO2RAbB0
siU7AzOGThJlbKNP0GHQVB1NsXG341qQV62KO3oDmp8VXbSs6KRgWxMzfoW/FGZ3
+lxHT5kWQQGJ8R2VcD0q2x3f1FPQ97fPNNX2fF26h7rllpxiTBpm3HfOW8L1wFdT
5NyiTiozWTrNTPEuolocQHWbflFzUnKqAFDuOrDxsc6wqRUKRZohgZU2TtqF/5QR
6ST/IW1FpKgNPGCzaERLFXWWxq7xhBvMTqt4zJ5FtHbg6UwNCKwsZXZJ/DweRk1e
uD0wMgunxWrWv7FzZcuP3GaljReCckCQNWRBlzAHczKPkTkctWAWPWxnUmG3Kk2F
jLu3bUwn2rzYiOmZdmLgalaA1g35jAeSUCZjacBgKMJ9bj1TB8gLmDPDJ+aGahyb
janbw09GfQzIck+Ptaq6BpBV1ZZd+E1eiIjSDxCkI3ybJPbGIi82M4cs35xT+qX4
skkgmUiU0VEMA0Fja+wGLWbAhWr2C6Tn55E0GIPrlUYlvTTCCPYwnDm36kBhONtD
2ZdDPo/ZtTg1sdH2xZh9hfJwjkZ3udMkKhzmalro1cUqK3xnM5HE8LV3F8+8zhg8
uJQaJr1bvkTu8pKpi862bKhrp2PpsutUob7LTf9PlrknpGN+uToKAoBh5ocilRQe
jYwRg/DcOhoBy8NcHGpnCWM3BggORsFlmGOyD/PgMidMhckRYo11IZZJs6EeB1p6
vJhVhXbH5Yz3i2GIGWr1HFUyITda4R2eIX6Jpuvm26ZXE3/Su/Svew+mR3gXRQdp
rx8LFKOeio9z3+FsQX8c43knFNArEi5Xgh990hxQw+R5m7Qpbld4X7ai0WyjJGFm
Teg1DmNB+6gSPdmlYyiBTJGNCNGxJyrYaf8VQfCy4V3KH52pawF8yNqxSmCoT15Z
JOSl577+PHIMGl1KacCPLnVkkapHdxr9IQWOihhOSgiaMbxzw9Z3+O7/IEgh4O/R
SL8SYsmLZQKRxthk/0AxNz1LFdBqVK/XzFUM05R8rTJ2AcBgcgaSEhHzSvoYWOcY
haKyjS0bv++oFU6ekJXwToLZr7LgMfv4V+A1eT5kjmUfsI36/5z+ZSPe4P7rIXBo
74JicZqklj5E1KRLjIhph0+YUs4mjqLn7TDhmYBobou/b6YKZkKPY5ulFA8Yfc3E
fkokkixQJXdRZdFO39p3TAie2FIAIURrfpc+IqT4xwuLM5dvBZ8SI5eDx9arhMmr
VL2Ylf5ZUucxC2lwmUFmZLmut9O9DogzqDqoDpMpkuhYCRNHO7FWTiKCvH0bdKD/
WRB6walwQOa9N6vY0wsFPEP0R3E9fxOIVb15lGVCrs6ymjndoN4qhMut8XcNE9f5
9dqgK9VFK9/Nm030vh3eN1KEfxKo2kjp5gU8B1w/I9HmGFXpAGfPJPIxSTeiuWcG
RqFG3fZ3GQ+ZWI/YS2Tu9bQwju+FTVg484MqwUSOKEFn8qzGJ0NbdVHtRKjOrwFG
yjVfmko7KEzFaturjjz7ommmv+hTYFTNu6eVx1GKmDvcmlPw8hF3MRaKPlU03vBk
Czfa7LR5kkzxLFibM2YQ6aWeqB4mjzHjidoyrQBHvyqn8B6XnRUN9PoWWbn8rPow
oXwCV/t5EatS9MkyLg/ju00x/gmZHOKsooTJMU+cDs+OcqkTjb/xEp7cnbxpQf6b
usPAWiJX6O90oJ8yYktwP/C3+zEkjffFJsi1t9wTBT3AzyDPFLbZPZKjJhnWpg13
HPsCLDCyq60k/sJ28t42ZOcUsLqMFw85HW657zBMRG/0E4NO734GSnGIPd9ZF+Yf
uRSNjLauhVpExeHcPdy5lwLW9A/3/DThq09IcMFzkfR5Fi0AvCDocVC9Ie1Duvy5
zQcx+cgeuXXOQvsuPpHhYjz4L9gv/1Xf+Sg+ejiXjRydOIubvqjmA/qw4/z3Emjm
Q2dSDucWCWzB7u0CD1f4/q2V6VmEvhrfyLFom5RQvAHaHjW+VQLHqphmT2xXLXGt
bjTGP8axRyvyPlEvlIBtkwwJqrV2vBxhxgWu55SgR15YOvNsnk3EW0+X6dmGMEDE
iRJAMNWF4ddGqqzBIP9Qus6c2lGuO0eitcfkrot8AqNsRSr1n2BnP9U7AfWTQYm2
sTvygtEfjVhovlJxYVsXx6WsvpjnNrcQBjedgW5rK/nHxaiFjVVgCprVKrGZYi85
r5FOVuCgJRWb9Zp9ASQHPTDd5BIc9KCVIt1Vg2P4CCt70D0pdKBY7DZYBcqAqJ2D
w90sPVs8n7WEL8ekcErYpKWUCVSItiFKf4P8s9E6r9aQzKbXoMJW1hHTtpeUFX2D
BCCIlQA4ECt4YN7+dC2H1FkouBg04M1lV7BWdx6MdS0NdMrdYSKYaBBOvujBSVF/
MqxX9xuIlJ9YJrahyqQdbsPtdQ1FERavTgg8zX0xhITGjK4kAw516T5XBM1LdODX
ZEc74nBCaSDlPoKVMUHGrY0WhtV0p3S9mk00j6dXXkpC2XNEZuVW0co40uu/rmXb
fpyQ6IrYPE/gvpEpKJRILK2bAAbb333nCT0XOFkxQhNZpY0Cbzag4BxFUF6OP9Vh
JE8y8E3kLogTxHDOFGdoqaYxNlZPMSR+DqkzrrmhLdq5Tz4sAyZVUg13kkvg0Vaw
blbhawE/MUnxM0WBm2RAnmyRgFTqEUg4SUNvX6hMoFsHrI6tqFW7a/sReNgvS0LW
0sXMEaW95NkLvpu/0DcXTyx+zGXY/+FDCBVu82vPNyoasn+lPNZFYrbA3qJcWyOe
vJGP5MDy5sBcLhiri4QSPHpCb57m9IItlvucMltoJ++4kOD/G3oOn71Oz2r5qNXJ
iyFMJotgPvalfGlF7i+f81ESrm5Ut95M4Myb1fvLMl5Tn5z02+T62SZVokQ6sAL+
XO99Lf70a+A9c9z8PaRicyLqs4c27oezyFVKJRGJs/4ukk5ZmXJuTIwIdeRneqZX
lrBrkIqLfVvVblyHHMyUv/shKEyLuqJ9j5h1FcHcjOqlYjnFJg06iM/4ZbZ76FKZ
V+rMfvxOqGc5U2O9BSN1FKYoMoKuAWqIpzW+WaFfzhc4VL73bWhOJ1iPDtwS3VUX
W3zOqbZ+VTbLHHxbw3PPE3Gjqe40VwaJ6gBWK0VN3gwiRjwLlxNtaY+1Mid3iIDN
QmAzlnwbf7kaXztqVmQDE3VSrDFg3zqgR2JH4ni3gH/gJ+X/0UWoO3WKL/71BkiX
4tenpUd4jay7O+1EQEISYnwaq1mXlahxWYSRvXWn5LESZheEVS2L/dE7/aoD6qq7
pn175fgvNsJsbAZnflbglyCXb3HYos+ijpK/FefvUav9EeDvbeoeBV939gjkekUU
W/8GNmgw4caj+NWYiPWLMB4G39LbQkIHuavS5iqqVgXGsA3CzpMuyXNBKQN7/teG
l2P1/tXOFO/FrnhV69+uw9MY2QiBqpW1VWYwMubzgZ0=
`pragma protect end_protected
