// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3x9C+cdtmKoh5gqRo1AK8q/OFEHFpTOVz08MKOYBjy56HAyVlqX9Z+yMXGLUJvDq
fjj4rMJ31/iGI9GBTlj+bO9EXJjhPb4HEI2yzfRLZE95g1e5BTFc+/VcF2yAw5jF
kSu4Urc1btXoYAaPJFjczL2cfjaygEiRBj5tQM80woxGaWom8DN/Xw==
//pragma protect end_key_block
//pragma protect digest_block
PWB3guE1glSobxoc5eIW6nmnaVg=
//pragma protect end_digest_block
//pragma protect data_block
RgJx2T4Os+QgEIRrAZJ3SKXBTnEu3Agb5nblqb+/xWPYugZmrEoM1kx8v3yXk4ZM
ZbEVdVDPhyj6l+jNkqOZmOdUwrtCzLglkX3AQ+/V0urWPBb5hRQBBanI7PQaWSq9
kXsz384xdsIvtELa7oxgwMnOUB8AsPVLZD300n3wq5J9L06pk5U5fzU9E45/drab
43Mm7x/yeBlxzPsqD2szXy2SNm6Z5iiBgjD8CX6wAU1AnOHcTWLcpdENvPbzAx+a
UXgGmlorRVzptboXZP0CLzQDuH2BDMFCuoerY+yGMW/3PkdOEiRsrdpI8/aggeuZ
GhOmhU38/UFLtIsi7QbjzkZzStuP1ExSKgglibzn9Z5zCl4J/vsoN9fYvZBmUgxu
DNMGCCjspbHhzyZWBhqPSPh9j1msDIxXw84azUnMaLyQGX+YqoIuzapWbveg9N6S
5PUZ/TRPMETMbmt3/r6ZiRKL5xdKiFx61gXR/QYEYdiuX39PxUHSsdEVcKwNASLS
nGlQnHoz/ilMwaRw2N2hPYzCZPvpr1nB7EzhbEtLiwdYNTGA8V+cI7VYS0YxAWMz
p2yo0zSHTmZ74AlJZJF0PyfLYs4KMfnJQEZ4DuGqhJtkJj5G907WYU0EPbggYIdH
ibElgJnkH0SaZgYTzo41tOBEImVlNxu4Ofspg+VljEsDfX9W2LizoVGQ4NpwKmYu
0LHKbcZNWiExr84i+ZvwE4WC/QZ4b6c7vnDzA1a+S56TBI3VKRX5QuGJRFzj/Wpc
LMOrGP0LdOc4uDdJSJpDQbzpvmSRkQgQsRYZ1PrlsqxWppzuk7Y/EvfuhxvSG9+6
SBdx95wkmObNKsAuGU8gHLp2Am7KMueMV68kDwcI13Jak/C8hWGUYvZGtjL0Pz2m
goKEU7Xoiyrun/h1/0X6LUmi6/AoImEf4KXMbCT/MJDIt25GC5RE6vNT8YnGLlOm
IVk68J8TCVGZzd63K21JVi6XqLtgTUZQ/CNj61k1BeWbGo3aaf+aS52TNxo72Fp6
vm+vh8/CUfQNKLKn6qjp6Z/zvCKaOl/Y0S/VVYRZfrreAyNOPFq8JmYbmlG+ebuQ
skhn4KcWv4+IyT4F31Uj1jMb+3U48p6dxogYFgIRhkFDQFhsAenSVHv31ZJoUa44
5J4AHSWhTpCnIefjISDecUCTht7D/lZ3tCYWXv9arNg0oEs3TzcN0Lf1E1hTKh/h
0l5rALqLicQO9/C137y6JLBHNHWBrrw54hGQ+6g29GadWsTOK4NGxkxNLwo0Vtzq
HK+F9qzKPELW8nfnhjw5RkUEa8aHvd2qk97Gea1iq6VauRdUokZQqoGxG3701oP/
BRUxaBDAYJIcdTfjQeZ6DTWUF/M9ny8ambHiL4CishdVxL8PS0dcVzMoDW3rvNuj
TKbf92IvsR8gdUKX/59AXMeS5fbEY/FAwh8yyhJHBLusLWqfC5l5Nm9B/IUWEvSI
MYiMy8rDG0SC4g7lpa5LHt9IZohfZdiUBvnY380DAN3McY2vukTU6kOmVZAAmV59
vfWzexxnmIZ+L2PdHx9zx+5q68AMYOQzt3dpclg9U01wwp9zV49DBU3qU+yQ7HNr
KfzcsQmOsR0GpIKtK9yJXhFMC9v8h80bGIy/WmIrsoFIYb/qHvCRbG4O2w0GUBV6
AQuV8mXcqOuHJfPARubB5Y1gLtJ2eKoBtv7FIR3aFMDtZrrOyhlqfZsct1nxm++5
voK+EN8upYxM/IZXdTuW7o2k3pr6K+ulV8qRzx1B2IOvc9RXtJff1ou6RlVH2vFh
G+cULsjaM3ecPI/slYXAlVV/hLOFHdGtalcJ111OkGsTG+2o4RO+8apjrL3ZSDSa
90ZEwEoBnG+1BrM/Nu5mGgK+7Uqkqp1T1jXGVx+LPZnVodbVjc1GhsKJSCCKDmmi
G7ZTk2W8n8GMbwN5qi4yAcz7R3qAPzcNh19IClCog8Ts4CmslkMTf/ZCih2oOvEY
bnR5mNrxl/nWnt5fQMqNzWailUvXh3lPZNmUaYn0qyuganPsJxpL6KVttE5TuLBp
U8lbwS9sT0eiJCOqYcCckBiTSCVEPYLmbZBkprO2SSXKW3aacvb50QKDMMuTNxG/
OnFnfk9aewW02SaAO/H9GElZZ1GExuRCq78nHwkIaQX9HZYNG3Uke215lZF9xUz5
1nXLe588XtTueSk2D9sgz4rvhIEiXtbweO6kadiw2yJMJlSFlshTqkxEqLMjNW3q
0g2a2H8ncrUGk7V5INmtJ4FRc6YJRiDnfKGqPqr3mmSy8XT9q1p9Oa/+j+Z2KP//
l4MFsCg/A2iYlmh3BFOx5RMbdRTgeM10SbcVUYVl6r78sJ9Fz+TVtx+hdOq7H+pD
wO0Z56ENJB1iFR6gSGN1sNnO6+pDHufbmrC+qTch4M6AFSP4CCBK4Fkb+ulZGkZH
76LwIpC9bIxZH609UkXZMhFMZ/6E9ugs4t5lBXewwMXQeqcTMEU5JAN+cnTuqprA
s6TC41qPBXI6G5MMY4wRZuIYgC/ZhXJOIaj/iyCjTZeKCoRhtK8ycJZWWQe+Nyrc
adE2f2bH8xSoSiO469rdwa7YYbYRs1ZFotobv2wzydxcFw5dFElZ8I7xOI+93JNk
RantA0bhbNkm2A9/zGVhjKANYw9AzY0iUfGQ/mfxKgs8lHVwKmyXhtuIOTZfaR4u
LCSDBN41tm+uq62EC0BA3tzbYvjPXcIIQZ+Zbp+OAMudtKlui6WaWLbpPUrKLT6a
hlEfQoC3qhTiLQU9MhNpJdOvrvixbMoMhY9fFHGkyKVOfAJeK6LQ1/ogEJYQnpg1
O1ZcTdw6B2GCJ/s4y8jgnBnfMLKti5A4WqCT54T4NCy8qjOwCuT1MgkCmf3nkfxU
b7WP68Y2sDeu4OYcsF0LnHd3qlQp/cbgGuar5bx/91DO/EPjhKRXV1dm2UIt3DcJ
D4TTampFTDywgd+F97fDdA0WQUHcSsA89wtjkUwHqQhBmNTtf85tjHllfJQGv/jm
0TJQuprBPJSEWoK1UBasGH3Z9N/NgxGjjVCono72EdnPRHwqpu5nCUSnckI78BY2
AjjGHpnHGgbp1Q7UE+zqJxubP5mVg53aRR/9nWd8rcvIV/dO2Ouki4kQJiodYQQt
bvyIPRLb9roFrDiOHTr0VS11xDNXoVuZePtI8rbr4F4eLdR0qmQPlpK/LbkzCgge
tA9vfAXXsiEvbFnE8kzERqCD500ASussL7JUpVsE+Ix/yUmgTgvzRYZDhvoWHLBK
IdAdRWwnBk9p1VYsc3hYdkHMxrdT3XdTyKx5/H8RUeIHliQjHA1+X/2nXPWFQ9KM
uRn2JOoNcMd4MQMRzBPxOnEubiHmzfg5KIzsszA5cx3r6G3IJIV7eVjwXxK6yMm6
7b8KbIb1hWxVbh/07n224V8il95jIo+mjF//SjbT/kBu+UtfrylTugy0TC+W+rMt
PLtIsqECPJn3Jqwn2Z+W2MLVfXDvWa/SqjXjTUZbqTYZL4xKhL3CCWsBjWr0UfGT
ThRCq1+y91rDYWKmAossYHZvC6EalH7MKjlc9oHdcxaePEePxgPFUzjbGAPmICAy
W+j+kUEPcWCxn7Kvzz+UyAZNSLewtOGj5WYHiE46TCi6ZeW24F6dFRWCxm60Q46J
GTklXnkXsZ3c9pRxajddLBsWBhgGq7InToJtDna1TEUrMN1RcNjOzgGBwJSCMJvv
HDV0ABrSNhaWnmOVQgoigqGNhfF0tYbt1+ZRfLCMaNNqhu4/6Wn/pLXcsWPhrcft
I4nXimO2McbaOE2r5VCI6FQfMdc+BRu1/Djgq0IFcC3oXOb86hcVJqu54mT9lVu+
nZxASyjwLDbooMTPwZjCcKohxoOMVulnmo85PytloXqUyK8ohUGNxy1F/NQp4i7B
BLjt0TNmu/AfTB059OwFC1FRMfnnqHXXEAgTcCgk8d0g+pcgf5pVF1/RUIfKT8D3
z37A3X4FQH63tO77IqOJlWO9IEKKEgkzui1Rm2TXa4rqtxhVHUO8BgegLKmbLOrs
Rz4pqohBxKCxj79U91LJTAw7Si5rhqABOWSanu8yuMzDQi/kPgSX07BA26eQByba
3S1IEkC8XhGjxxxQR72bFpT2birHuT5IRH3TDMcDvfDLlo82X9ovhDimYRNj3/xZ
UPLbV3jgzS7v8Ui9g3g1qBqV9aYAZksqXW+MKiEaMFHq/L+4d4rjNsH6Y+DgRHCQ
jxe3lcsYB0SS3BtgVMqCc5gk9V1rHZAPEqNufQ5eESLIeIY95JdEHiYs811Pr1qQ
T9CSi9SzZOEJ2Vff0M74bXhyw+knZurtFx4o5dlkQkBWj5ENtu5s7pEJz+eRKYeI
huLBAc/US0j0J4P/hAmfWatKgu6DVusuY5AfLF79ewr2HgwAIfbPCQdiKkOGhZWi
KaL8/VUnwFMbqUEnf/Wc2AckpFvrADJggiOqQ1UOZwBc8i3i5wCo6Cd33FMbyudi
rUqnQ+Zvpfo6+ajYfbG+qlKIHUYsgEQYPqicp/P3rdKyl0IBHsRZNZluRNy/7/8O
dCgrbhHXJPqlvtDlpRIYrW2SifKwHwcnEpDiELii42PxkqdL8YCtmiSWdacuU6k3
mS5Hn4UDwHXuM9g8zsRni670xwnE8rlli45Xwe4kaIpWDuAuweqQQc15NzuD6G1r
e93UVrGePhyfwN0J9akFwTfpabWrW6r5KRLudQ31y0tfZboBPEk2uHoWJTUll9ud
4tuNNUKZc/qZb10A7mZWNAZqFU/inJhbdR193NTQlH46weMl48O603NMN7m+MWsc
an2bwA16F2Ivm8ytDjKfcbcJgxN7gDwOICD6yeQEdU6md9DKSDwDSc3OS1GhqrNp
v2NsQWKpUM5x4JOpDDy9kvD1SjdiRvZcZheqyJXiyHGwam14+L173aLk9LX17XKI
v2EQ6eesrGwyX1jI3PzSglq/4jh1fEEhMEo7lSlSI3e3CXNgPXJ3e7lRKAvqdCVh
PmzKI3ynDzU3Ljqfdaklf/AAGg5bTc1TH9aYEXUXC1iUjdmJbhj/gY/7zTFHncpL
ScoqT1r7c6Sk/5Cwz28KtwgJV5GMc5S4SShXTKnuCcJ8naOjONXmjOnICYfxWpAG
oj43f8LXfbVwOjirkSQQ1rOXUerWiW5L83TTUi9u+AywWOaom+j+YzWMJ1I/2Gcb
HAlZYho8oAqF+WgeNkKk+WprxV5Q7Y+5npw86jK4N+Xtpch1/3enfjCN3u34cW6E
YDT+1Lmuf25M0+UeON5aUtYTQbT0FYaZBYjQD4u5kd7KovDtjhBcWdQizB6DhY1E
EjuiJXCl9VhTonA5igs8MQ3GHqBiyYzfrTUCpMWrTd7GaF4RCxGKijVRp60HBuhP
yYWBvy5Leg04bAED4peEA3KpqbHp8xNl77QnpbJZjS5g1mKfNwQWT+fItHIvqMtU
KPVnmHfb6OD2rHNhn3iOV2SE5Uz4UR9F5dnvjf85u1K5K8mqlQat0U7F6IEb+u4d
iyqwDDAhfc2a7fDLK8eVbwtWiXKW3P9nbcSMUC3PHFoJvITNot3Wl3ioOSIwrnmo
XuArnJFWb0Ryo2+6LXaxRxDQp54t3HRAjli4Fm0sWSVPDb/vR9HwMERnPqbrtXAk
R9tynI1uENhmHmVRbpfN8x95NOFkUBMtX3gJhyloTWEpHQ4UoU/zIOF+F+lxi2Ex
mlCv/IPOwVCGzbzBAVNhHe9UCy41/isZetAFZ6Ra/t/AuWIo9qwQVpnubWjRL4UE
pgWMEj8B8j9Tj0I5bTM46hFni61Fci74Xy3ZL8Zol5PG53h6Du8vuOo37Vlx/kYX
8bBlmFh9Uu9zNFKOH2V4RFbgN5xwYqqoZphWx2UD4TmCnDRUQOW/QHKFV2e6bORC
/2xcWcNqKabycuFHlzB9fuaVtXVvJrV4NE5sTcr9Unwd0GLX3MsDkZoTG76imiYA
DlJW7GjmtqWXFjYt1OmUDIb9o3feh01nR/CB7IUF49vSQRMofTOXg/MI3KdgTHOJ
LpN6G0tGk90MUrWLNAGKVLEazYsfHxzxZbmXf3t1WHOFb6mqTssBw4muk/p5r6HF
n7l+R+/6ITFJf9xQz+g7fJjhXXY+48h96IxHEDbxObETpyBKcuan8JNEtHv40uzW
bM8THU8FCX+CwQ1jmxMHvHhlobVObnU0Ysq4bvB48Us16gXJpCWFRsdEfpns/yI0
sbKT45ZRndcLmEvjdbN5a9TTLGrM6/qaZdi2ro3USiuQslAEll4ReemkmBgbEpv6
3zmIDA3ULhkhefSpRce6VhXmHYchHOLp+cwsUlNjWsG7td/adUP8TYMGJJApoG1w
XgM8YrSshn7NeInzaCSmmFF1ZPXMJ+CFPaXZB56w2KChda96Niw0bDSfSLq620tQ
JqsGMuBcQ9xbICasCBJ1yHRUPPedqimvpwE/AX6OLgqbBECWkYV8EhW9l7hZ+Hf4
Y2/uNIgzzp6fyHu7KPiF1Gfr+YxlSx26GxmSFcCrfUR8CqqYpRKAG45+kFpQ0BDM
Q5iwb81HPvS3HEg+8RrDTn3UpVFxyDCMrk7pI81jyYjCW9SUHHees1Sml1vDjfr0
hrajYxsrzZJwadj/Nk7/DHg44eXfGkqhYnYpxaCU4g9+ZwjJFMUYZzPrFPOEO3wl
R9paY51niX++L2WbXsuOFEiqJRBxUpEsVzymxnovX9mSsc8e6FSgS5qDHEflIkQK
fDsM/c6X7RrD0R+pg1SLRrWxz0K5FCMMF9jhPfGMt/qg9vUAoB/csPAugDZKFnMg
NU4zGcltaFLmXc8p87b1sgfidmovEW5ug4gbTwDdqHIm+ALQ026D7uKUHKzo33m8
hMR5fCx4EI/UxypnBXtxgec4KXjPAKbxyKj0P0s7CXG8Epc++2eKUQ000oWkYrnP
ewdXyz5FrgykI4AAShlVU65hK21xYBcwh4WEORdWsHjWg/Gk1GB6Ds4EL6PsAFL2
VO/yvfDFTuudgSNtM3prAYN3o4mgL1it7SZQ44xkq4zhgnNvCpNEAedZYUHaBaDB
fJGYwabYffMQdnrMEU7EXc/dbv/Gt1BuSF7Pw/3X0nJvI4wgqL3NJN5UOuTNmVjr
OYBGrO+S1TDUrSySntwFlGnUCdBOgSq5SBtcl9oxysy1OVq8CJMESxqx3ApWNy7x
bvXD5xvQsdGlI9uTNiDZlI5pvqBWEjcnAmGweF/9tPnfycPif6jDrDop22NhbbNh
cIAWhnrpj+QOtwwy2ZlBuJ2AP5gPkr6n+tjqH+loiIqew59u3MJQAP/nZ1CA4v61
9Y8VoY9450Gbc10hHScfGvladU5HZap9+XApifFVE4/XNBLb0Fem6BYHYUp9TTgg
IJBQFRN62r/EQ0I/kEQXqjBWSmIhtCQ5fnoPV7jtsO6X+vQlhi0eeti6/pqVQ0kx
PfBJ+tIinV1mIWK4vrW9Nzagf3viwtbPXKK9hhqjsjeqBJHbtIqXZyjMgGLK2Mpv
j0gwINSO6bGCZFZp4u0Cboa1IX88ULSXF0FiiN867WblNHLJ461ujBxKhCFXHhXB
wVFMNPhFCXniR+p46vRFPouDx4ZiNNxxPpcY2BfmvKEI0i3v4wFtHOiqs08KCExC
+CAk88k9cfUbMo5gtQY0zrZwkcBjEDCbmC/WyT4oozD7HhOhCrhiz1o1tr9iLbm/
Zx6LRNEmYAlW2uVZfmcwU6nVduHqnAeX+2x3Spc2V+uIg27D39mUG/tVLgqSUjWY
zNBS8PbtxCcT0dtoecbvRS9454Jczcc4IJ2G+TQx3zqBYkVQilr5qJP2cAo2grIH
pIRvTuO+Xo//WRdc6oNG1rHw5IUFcUKwgiPVT/2tiuTROHNpLQJXYZN5u4f3Vhbm
mw90h6SJ4zzubHQa3in5NMosa5DZvehrt7m9FYNiBNQCOVgNxrjsedeWC1oQioHD
d2TlwzvlUpDt3D7c0j8Q3/5DxyclJknn6z8kOVi4Rt/NaLydxB1QTQWFEq17qwR9
4YybNPoGy0rukfuxnC1g5+ghgmJWXYYI/z6Ou+t2n5KnujFDyFIbR69hj63nzADM
IpNF8x1LwfaSXPY1SSqYcuc5dCU6neA+ibRCPCHI4/LnImKPPzjOjxfZIB+Q7/wl
wCUw9CSMX2TkufSIxzEQBhFQLhtqfnae3UfAHhu7d5IKNSx2YotaF4/2/nULWrZy
YTDysV0yvMIiv+W0thLHRIczXC7E1XibPHeCvrJ2prbMfpVbPTNbJs7tMLl+G1ag
iVy8VT6pijYl8CqVJo+IIiBlNeB5uF1irJ0I3PvFoiSrV/f7C3hbGRbim/BwB0E9
TUAY0FV4CqLzbFu5+ru2ybptyJQzG7wXXLZoOGeB+pSVnlbstbkrC8pMUN18YObN
sEatBL6pBcvq5BeMTs7YiGCCj3XzyACnPpj8hViVN1JvXeXczY8VtwgFGl92GM1E
WpYIV7swc1HlskXcDbskDPRvlIvSPxLuQemb+EMY9NpNA7SEzFQRqfFpiB0Q9MKI
GCGS7Kz9WrRDElkyu5uDXZ/P8Hah8o0HQtFx+YBJ9YzAD4NcUw8UipFCjxtC+EEB
iggNxTirlgWu/aaiw6vsdgQsFH/FapPBrEUiN9Gt6pTVR2aArCYb8f34NMrXQ29U
K6xnfASenUU8HliN2a9l0Qvv+ZPKuYjQJdJ6ttv0XaWviy58mqWyG1Mn2YFWp9hD
S9+XoIGLULGvhyTyW97zBm267IevS/oVS+owiAjvKGcrvvA5QA7HvgARqwb4udEM
AM2A5eGZ5TIZPyjbliXL57xdt8ISQXEfkGASOH0kqz+Z1jbHhlUEtyWqjQEEikjk
2AECiEY9Sx5F+7CQCFP2hVdvAnJMSSHRFmhlm3Fg3he5EQ+li2IeAxKY3q78qsWi
5cEm3+bUAyJ8pRpCdEAoblrbAdj6DzT4MeMeIV7Or/8ikFAk/u9WjqSLJCBZ7OIQ
/QSkxvEHTEL2zT2ahYmBSSbvAvNLWbiBaG2x85ChQdPktZXqKDpFRnkZ5ktb52nG
e7wd3n6MSn+CboJ8zRv8mZzLxZ4hf0+dt1GgGc7RaihWMpTGxsX15QxgGC88Svbj
KIrZXevSxE2wxxRRurRZqT/hVGWZWhWanPHfrpKjms849iAyclw3iyIb+XY8H+tk
rUapZKcEXsT9lHt9DFiMPjAxO/QbRkYWTMuR2Kwc9Hkvw9HvMoE2+BO/7C5RoEXu
rsPrDe0TjUmxmM+XjPOLVkJyJ3gi6KWfuNi3f7GBMx9D3oQsMG3UyG9Xz5w3AoAl
Zwxf48G152lwB/rZwVqj9bJdBzh5OYIExmr8wYbifPmGYynOivhtPsB9l5rDfdJ0
4EjfSTdQWoVeAaEDCK4yMlAgMNv74pVCCEbkJGT9DCmxdfZMOXCf78b+AZlDINvz
CqCMMm4f4fg7Mj1zKPqhHqWKtbvj/8A3dYUWIJxpLWQij+DfNNoBKpR6IoIO/lss
DTUcQJxGD9cfHqFH+BfQ7nir+hFuZRFCyPX8gbC85DUPWP6kW6t8KmYDVQoXuURM
hz+14gEeP0VIx5DUV33rC9rrnAUeOwun0N2RlEcNH0yd2CaUbmsbEFbpggZ4EHnT
nAyBXAftwTr57DMRtCUEDBNYdDzr34EQtKs0cu/uH9jIAkVK+0ZZgbWiotBKmL7+
IWdUH6uvhDvPGUg9X+LpIybLohHSDrnGGJ66+q3Hu9wldqlYFKSoE86PprzHnnSA
AP05Zn8+no4V1F7gRYgCH3iRj3csqxHYiGHQ2Q85UzCd1Ykye1LB+kH+krzczkSH
LtHmXsPXfsVqa451AzOBNPmCYHiof2VWMQrhZukMHS1SGvlT5jj1vp4V8fLNXsee
fLMdiCUr/6e4kByIfSjwWsYUVQJhOdbD8EYi93Ckg2WWe1EsqNvWrrgWMivB6Azk
KSqA69aVtjYt8qtGs9dufdMjmZeW1GdzEazYsEmokwV9P1D5NeoRdy0gMscCEzoX
aspCiJL7xyG2k4YtXzljypiATooRv6d6Mk/LpnXRpP3Y6gp7wduGdtEYntJrs9ld
Ue30p32Yf5rcnSLO2JA7Tztl+P2TZPIg90HvVoAGRNNJx8seBJ8JDA0B6TZzvFSw
QJKxqEBacpfxCZkoKFy18U2NpjlPHCL8ZT7PY6hn03RlRpLqoJkRSp7gnjfQwfXa
E2umw9QvJKbXGcX2XouBwmFsVl5/VmqDshFIhAJDVTc9IsgPFL/5IHOgoVMUnUf3
P1pZLnk3XJ9q0WqfBwb3V/pd6+WpsAPlc3eurk76Iro1ASaGQBTsK/6PBnxwMkdZ
wf1/rRK4dxh4gjPYOvT7tNfsgiCfW2pDvAcdsuc+ROk8oZpzfeH71A14QRCMCd+x
NHiv9yWrG5OajoLpNrN83ml6QkGI7tt/jhMDaCd5VZzecoeU0IThkP7rfR0CgVVt
XnQ7kPH+tqvye1EW4jhH52QeAHS2l78tVzw0FY4N+pUL8NNV0h0FZq6UeUeO1CvQ
tHsnz6Zv2INcknLMsOH5wAtkg7OguHbA8/20QSJvvXFkGfJVwfGt4k+MkXHEIRVI
1h5b/66gkw5Kgimwez6z+2extEIrDUY70Mlvdch+ebc/HWC907ezi3GyhTgK74en
0cQBGtrsYx45TK2MQw41lKqu+vGFFTK92V039Oy91aNapdfKQnU3AdZ9kiGvQZrV
LzkMSk1c3GFkhJZnLWcUDBoEF4tsMm+/HaLmKTbWaw9uC4XIiWRQgKC4npml5T1A
3EFioHZ409byvYCDh6crOabqQnipWf5V9ezK2se1kGHC+GcnQ5WT58IYM0qJvF/v
XG3z5pzTx1CCVrogbVcmGLPRDgkMrZuXU3W0bWeuZDLEb7qPzWRRM1Zf1ElkUx8e
RUwXYOildDyo3t2q6fEAnxtxGQfUBTrPUMaGhpCHWTQlbvqEptrneL3eulE3lB62
EtOWr4jJfZQsdAapMjIo9/nPIhTNOL6620XBCiBZAzDpjkk8vdvEvoeOX0b0SCi5
zHcbYX9Vu7eXof9GIZk++g2nKsP0SeBUN5k/TNrfq7UD5stn/BJ4Lp/RNC9/+Z2v
CuEY1EUzoSlmVxwwmLBNPweNZ9YhUucxaI+AupSrAoo9y+H3oNNj40J5A6Oz0dRD
HpuUa+4XGAfLuHDkfufFMaC1OjJonqajeCfzP6X0N9au/XjBPv8tbcP77R3FZBUW
i2u5W7bMh3MIGDZhIzBChQwoErnjfzlu49aTR9/oH4flH72aJTIBljjU47HAt0tU
CDez8RdUUfsYotN4h4mBvizFOOvWWLmmYW/WLyW6AX7YFG7i/4tgtP1LxLyaqEUa
nyp9nsAIDrMJAD9Eoix5VTnnXedVnYCYabytHzwOcQ/NHJwa7wD5+RxUh5FuX1Ma
r16TgTEgQsNe/c4a+GcJalmwATJrl99HNOCuRDVK9ecdnjIm8WGd0q57kzb5rlAs
bmKA8vxcNAkXmbIqoCvR72SDrHeJD873gH8AsW+hRP452wvS1ml3neVnirzySiBb
Afu7IjayvFSFP6mKzN50UN1jLZJt5q+XTcJn5RC5kNvTqiJ5Iy4mbAYNZyvFL3kk
iD9UYhLwOEtdHrVqYF2qW1iyf3e22UZ3L6P5YIyJLyX24zNOu2j336Bn/i6d2E3K
gceveiKV6zK993/8R3mlOLB8ECdZxyd2/qPzxGSbHR2dLjm7EHp4XK/cb75/8Z+y
gpCEbqgTsiAsCWK54kH9nsr49L0l/SniReHIaCQ9CtOpfdaeC8anQ8gyhHp9GEKI
rMsq050DDAHaxnP4H01tVJckmeXTksZndyHm+MmSdl+pHtm18hI46ViRaePqpbby
Yyq5oPBg6XdLLsybOsyAVd3joc4d4mUi4U8yJlaITxonSFPWKZ1GAQ5q79ncngrt
IGUTlF+opMfkzM+P/GdrGL0b7Nohw+nSM+rn9uqqer+Bgyt4lg382NeAK5K8pe+0
MonTGDjmPzTZI17IkwPc8/o2Y4A+CYd2Xpt7yVsYUoBa6fPhmWDhVnJciGBAOKBg
VJJ53y0e4TYb45oiq/wnHFmZ5mSB+b61zeu0ghjwW/aYtvEXjwP13pr1r54E4jdH
5CtmSiC9yaxoVrZQqzCSlm85eheq9Hysgho5zJHdXZlAH6RRMzsatTjDLnIPtkaw
+Hgg4c29NCwr+bLiF5RKJHGHPFaYYLeHvqJbyTV3y8wFeTZdUhrLbbbZvVCVI94n
fns9By//g6O2avF6xyOtJ40s0upXQMWHLYSDRBmZ2AJFYp6z+YXzIYvPQWUu5TU7
wDJ4nEChrinFoet+WBQKTXUj+aEtId9wTMEIWGk8dvNSxkTLAfapKNu0Se4XM4rR
pAIkhwCH4saF7Pb0EC8NtwA0iVq93KGcGLNYxRjrmiwOoXMcs1ZF/VfGohPzfjjY
a0rXy0bpUJCKFJVgr3XMLsqaIdQGPsV1gPDsPHyLF3/Q5KV/lAtsxjKW5WSZeouL
GsINqh8BpD46RdtM6nBZg9ioYB63aJpTtADbuyQwuQ2DjpzGdKH3EeFYQx2yQ/G7
gnww+MnJiRQX1+hEEMWzHr/AMe2ef7QW3RUe/9NRnhKy0y+GL4OFKMwT5LARl7Vl
BiKDBnR1sC8j4pD394FTwj4RNo67LCj+5rGC0pAoexNdezxGYuy4Re5W6u+Kayhg
Y0q9Duy6NKqxzdtsUTIEMAQ/6VwIFlLrzn/bT0fko2eohFXpgwxX8nXHvO5ZUWpl
FTjbwwP30NuanyowTgbZ5mgJa+qlLOP5457UAy5sXIDbfQEJG1k8NfSD+xUex34i
lqKY5B7FTe8zk+ClZe+G28QRtMVX+j6esk69l4qPYb9espdDbKw/Gy/IPGz5nJyX
UBZyhlM0CBhiNuArQKlV6ICRpFdvGasnt0plHAKJrlRGM9ey8+DLaf/NOWvEq6T6
7qXu+GbAbp2sX6Aez8EAN/3mNC2/1Eyn5Q+Q0CdnXhSuBOJKoPn09gDgURxPb7Z3
w/FGlPhn1WfNYXq9fHhANWS2KhE4zQb9/0szrpknpTd2FixKfj98BgXYP1OFho3Y
Rf72A2NKNN/3FcEZh28NxXUzXRKwP1k2+cay1xnWWP6Hc/pYBBxP/zKKq3e4BpjB
g9PFFateShLWJd3hyTbCnFP5UfdUqWkNeZQ+pk9R7+V9dwNeBsYBKLIXL1vFIoKv
9kzicL463ri0kZrVqdVyEy/eexCR6x/ss9Dlm/nc0+rSyw+5d1J4qpeUb/I9nOqD
3Cj1xyRQLYkvgxCwiE1R3fRAfvoBJR2fL1TwjJgWHJ+SMTsfU/u4PZ6MlcjANyCj
QK4QiQRovDAt48WyOwXwovz8MRIa2LJbQFrCNTIWD8PWk7hoC74BtBNIEezu0xUj
Clwb+Wbe9Adn9oJM66AGz9tZxip/gF1UBV+FdW1rlAlIqj0667bxMA4LxIDMd2WJ
6wgzxI34VgsfQ+4BZEyktvL9+n8q/fvl3xMqpm/kS5Y1LZg7HLn+Ax0+Yg9JynvN
DfduRAA51tyqpNoH8u/6fUfGl9049RarzDf30tQWQJklThZ9vdOrptkW2jYqShP7
OSNn82PNw6iyj/DvBRQeL2ruLjnJDz+xp3gsh7vdJSec/xHhjlQfL0fzls6Sy1ng
g2WwqVEzLcBdcgtIIuZ0DrgTQephorvdgDjdzTmiNlZfiX7YL+QXUTGluGx6qish
HyAxGM270VnOLiaQE/iSGeRJaOOO6iQrJJBDq/tXbHZ6tqI1kLCqbz70SSr6xPsw
0j4BF22FT/yPmox5oj4jvYPbzoyQ3N3O0tlJlCJ+nfjl0KmeBbZFcUIRmtSzkeZH
mVuTlSibSkra1STqveqdtRnfHsfC94OOfOI3j3rlmlHgOE7BhrakX4VmyDLi5wRk
nz4DtG5T8Dda8TcUeK3ent1vggnD55EjlweI069QU/KOU8S2VJcpTh4Y48aZrIB7
J8IXrb1iFm37Xa7edDvLp65F2oCFuV5BTOT9XsWb4Pqp3qKkw8FXAJ+FY531Nnwb
YLW/44RkTRDNr+NrCDXmmY+BBzN9NXhQ+rGSpE1fs4srLKaT5wvDTKZ94MX0aCdf
J09VbmXBqCrbl3Fhrl7zYKVGwI132nHLyed+mKmLcn2DPy1TKAkilaZek0z/Uo+A
wQF1k6RhikuxepJogbqJ1zv1XNDytgp20wORpRQL+FvHCs4gJa/i3e5FJtz7MixH
9wts4DVYJFgi/ELMryOxsn5LuEfUCFhaLoHsK0pY9IavtBIcYIGlODmUBHwRzqSU
hL2T1nX+iBp3vUG58KmzfsphBMmVVlnDzuLrtfnbMYtuBlsYnBiFUeLlTpARPovs
RQAd1ouAT5lWB9ntiri0FMGCHUZLEwLaOZiguYfK77zPhZmRSnOp7Q87iGIZXSiQ
47CGTKbWgT4YtYarZOVRaY2ZqbWNs9gB/z7HLAOCXpIHwumowbtU6zStlNr+xy4A
TUAk5tkRmGQpuX1nwUDcNU0vuQtGdHofEKvCLp/HYZEVYYBg4W2sQEGv6drDrl1i
yeWwWysBL46EG9/o811/CoPNo+SCAPnyAQO34BUEXridtyozltcYE46qGd13I5RW
hAlXxEbcf17YtF4ctoKpCyJU8WNPVnL6xc7k8QRmh8Y1uk7p4mDuK0S5wORIDjpX
fw8aXnJ1cvU2+cI7P32NHQernH7i/Klx5ZKjMvH/Gc9ApH7I/V9hjyA8nagH4p3i
Rl6vcpOaGrUrER5fEXKoK9L61LWO1sG6zloklLv2tKmyu1IWsAfYRhjyOR/gAHJl
Ron14x7EZ+crSniVW5D5QNaD97dcs7+J1FlFR+/6lISzFkxmA2eUSIBFOdFGuq7x
ZDiku1do8kACV/bS7LpJpl3UEPukeREKqFAxFGgQ5x3bYqoZUMihQDDwKiEikWdc
xntAxNXqyiu6ry5Bhw+gwMgtk6VgtXdSXMhdfycSHXlqqLhNFV1/grDOw1pjU86c
a+zUP+nFdRrCU8u0ThKsQDEbiuwLjiYdLX2rHuTK9hUWqhkr1fm0KBYLQP89J4Yr
6ThTmkdXKMDdYP8mpde/LctQ1/VrH6iZRZFOYK0obpgdQfnfV5EZa7F9BCngVdYU
z5xwz4PUDIv1hkkV8NBvJ87lI/e8jA/b64472BDKPU7y9EYS5KRxkPD7G4X/Wqar
1U/ehyAtX0Z39VJjV8P0YaR/UOVjjE1VGSAZK9uM1cyBaRaOWGJcK1W3tZE0M47U
dO6dh9vYkT/RGL4Gc1SeSOzNe9AlJ8Fi2e1swaJjCUvdKIU6SFzwwZI4EY9SJJca
fES7cjvpvU+BDg61zvmrISOaX5DVP8mdyZgxBLkDnOcKoSd1FzAnmOKREeQSkKrx
LYD5mcQpmdp9koGCc4nEDF8GvUedibn9YMNuVXPNERMoLQmCB3/G+tvjsSXRXvKO
kbgTZCeDO0RS1pmhnEM+fTClSSuaKMrX8q6FrKBH0ToudCoDVqW+2Tar1it6IluH
yPLSvn/qyxxKiokapFclSpG+1IEiky4AxLQwBhyz43m8vlDwoJrQ1ww9KMFRUAdU
F+lL4VWU9MNR5d50htGqw/bgm8w3zghZoulNx0G+iCv9G5k6CuQjIXVx/rgxEU2Q
tmM3Tdpe9IDIj0xUPG5Fyr1GoeLH3jdCKktm+rUhT1vcLbI0TfAGNB51SquTx6zW
Q7fsCbS+0WiQNXLeZ9HP811v7hAK8Rt5Quq8KnFM693AjQ+R7LLfU9GMeEpRFFod
VZMcH1lfRu0Vi/YK+WmTrGjbQfwqAa52dWWcptU4c6XmvBv4PTHAEIHNiWbMFNee
Dn1tE/mD+vr3xctLYtBoN4nYUkGNTLq2oHvdajzqom5tlPCW8USUadvcmMyqws4E
CpOi35HQ8uiraKzapBlKVwovz6g8DFQYTuBhZT9HuBFBCqJRRCKMabjknwxWi7T6
TDtAQUJFKN3+fP6bA89wv/f3B2gWuQCCWffH9ZkBBz+pAY9CHSeaE583OPrNLBNw
10X/GJOpK48JcitQyLt0xWmM//Ltm4m4LeXSPxWAl7jipIEYme84j8OawAXHW6U3
L4Iyt4QhebTTlnysdHvGe9z6RagFuY2qfQKpODiy4yCtf/zMxGT5XQ3+hgF/tVg5
P6l7jz9e9P1kPJSp28TQggdIndALgvsq8GVGGuCXbRn7hpORgDFAvSwJfRIljkfJ
aatUuCHY5Bf1VRtk4a1KaOSQPSdGj7NbAP7RDRkwxCKiv0EKDnddvPksSDnfCC76
zpSccG+w6yjPra5ZzKw6avNefGSVbTkbxbRA2LaHBkH69d1C+eX4s0J2EVit6jRC

//pragma protect end_data_block
//pragma protect digest_block
a1TEusZLqSc0BOCfU6KyYUIepVs=
//pragma protect end_digest_block
//pragma protect end_protected
