// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HKAwlAiXrkITXQNQq0UsJpcMLdUWcL7KFw3Syqq32tvptDUuL1fVdyRLCa9h/cljDCPvgO7XjsTn
7/nfsh8us+cj5ilJbAAbL4cOzbXrPHCJYg4UlMBIOVBaQ9YPvksPLBV4zls2Agt2mItO6RjKDVmJ
53UodvMncB7m02PfDrRGQwqkOpyYsPkWUsKTkakB1ZOqSJ3xNaCGezqqfyRyjbiU+ohJVNno9m2J
+WipdVcHq99txdjX/O1aSiBvOKpvCQLX2J3qUnUN/yfuT5r4UdNhoi+bt9euo08ieqv1+bNPDffP
/eR78hfvHnf+HL+aM+UiIsduKLILq+F52dT0vQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
H1PyHPDoo9fhdehLfiab+Wl9M9r/hSseVjx8GadOS/JKm76XpgHvV5ES3domXaHwLOnTrEcWS+pW
/dWbSct+iOas1cxdR8OidIiNO/6nvWjrLJPtVJUfMb/znni1GVmMxa4yKhSph310sp18cVKGUZUQ
uzc488i5CsWcgB/VoYsFS1C2wAjnNE5zw49u1wGqGOkCgCHfCCCev26brk9wvXW0GsaEqr5oAZxJ
frmRbHiGf/LcCqdgF2YV2MJXJr3MAUlyhOnpqeQHsSH4/2NjsSPWMvfa180g4MyMO0Tg1sgYAgh2
jKvIWz6w/zYjWr8lB0jG6oBKolbusGAewEeuNXtgUsMD1c2T4OMAL1Bprh0c0c9/knSZUxkv0iF+
zBTywnrn3oC3Vr4Y9WGY+QEhDQyewCUY7kTem9/va8aU40MZ8tUyFICb4OZsXLntWJjXTJ2HL7ZW
J7jYYGxfrMYlkGq0J8LoUkgrNtotO+dY0KhmiiGIdZEp6CAI7gvWjTu+rJXkXuLR2OabinBDMOJ8
06WR2xq41lc8VJysJbwLBh+nd2n7bIpjnJMsOh4UgIVrGIr3mWyO3403kJdBmt714yuV4ZOcB2yp
mXiKlz5MUNwoFfiXRk96GY7f68/89BWxj+3cj0BtNUXSSK9zc7zWLDmWKeUsaRc+CWahtwW3Lx8n
eud6nnjhqnO+VuCF5gmT3HqYToQN2PUyPVch2Q4GZIALwV7lVKsmh18cScH4AnFMaHR1bjPRgRWb
wiDR6tcMc+Qi3KMQzcNi3/lHvNuRCnLR2zyLpVZk1fJ5EqERv/cqWYba3rnaif/a4SwQAc9dxvBa
/Nz4BX2PnxAKHGEZimLYwM8FWNg2suSYmTpGHuEMi2RZCOPjkPmhO180oJd1t4dzd6Jl1AP3+FwU
NhiR0OndaYNlEfY0uJyCF3dNnsVk8DDnZCyTBDScUnVOVR5Hv6KsNJmvUyYDRgKvK4hcKeRLiOn+
gTycuAUXEku94NBnaBc1wFdFE37dCSZLsGZ+A3cq609PA/G/f6wQyaQfTx2ufzggZ0wFzo+b+HPL
/62iFcmNrU1j/vNmaiBZqr0C0nV76lhSYxVlqGFriIoTEx8kwFK5F5gL0IYlAU+8cd6l902WX4/E
fBTovQnlgkFzsB9XyLcTt9rRgb4YU15l7nDi48X2o3ExGK9wXqvrQSf58KIUdnIrsSvJOT+6Rs5e
44+tl57YvUTu7cBudHWlpT0R6jzC5cykKcgIKNRyTq46lU7bMeLtgfZmskBP+UNmMP5EOATCDCyB
DZ/odzKAnpTynB1P2XVaGoJMZlEJXp2Gex9YEkOZmVJh1iENt5zVY2gyLkN8H9kYmf28pYwf2i3u
NETokBrvGojDSQdjNVIuaFSeG9Tdg2EfHtJVYcu34YFDzCFgY+aNGG0SCVzfSnVj3q2OFabaFYC5
zeF5Er2je2OeZti67OzsNwT9kLhbgApxYWJGk6ipAUJ84UI/0WsL7z4EXPVsWEucgQFcdpUCfbSt
knGIw1a+6T3n4khrs9Ojc3B/Pcz7tPJRob6ttukmH3EnNz9JvLyyyW1ZP2eBZ3S2Ib4lP/yUQpAl
+DqV8qsILwaBZD1KehaM9lgxUZrSlSq4IkVPuh88FuyExLJ3vb05nBaIzdt0yqMIFbfznumj5JXb
v3Jp++A6gN/EVAVI1FbIonr7Mj7sGNM5OBg1KnBQCAtXC9wxeGREJWEWe82+/oXMQCUpmymPlVZb
qv1w7jzfls1VlRvPcx12ymqGnEm7rglvTB5nlcMdhrrpwD3PHTDXWStJ2EEFygn2FYWwkxgfMk1T
LBwWM+1uCO89sx4ySuXQfAiWi/Qn3rEYOp/9o3Oqd4mD1cFe1fa+dieUzHBjvnProElHGPeqVZmy
At80SZ9EfAWxQg840nJJ+PEJeVaTQXbpsyws9DhN/cTRmXxYhLtNW4c86T3n9JR0VNR9LbEH+wP2
TKUHOEM66zw5f79ZI5hp+gKtKEamVEUFZ2FBbwZIY9MCF0/RZUM0jMf0rUNF8SQwrIFiXxHUimGE
o5WYfiMvczBm1ui8352HBDQFxPeGkvVTAgsk1AbqzSVkHPBE+vLsYKOMXIHEuNY7kRSIs4JBylZQ
4Ml1CJnn/MtLOWOyciaWOxjc9co7/jH5DXJK2ZqqZE8koq5jJfE0Y5PiRQ4UWQzHsHGTnLBbbpIv
H9kmYUUCPRF+N3+8lnVQ/UN3eIPK6eVVPqXXNW/8nLJNCiqzMWT7uTMzTv2mDxjAPDfQFp4mmvrb
4loGDmvUlbasbivxvOvYvLoOG1eyhjM8MN58VrTf3ySA7AU83oI/ZpiYX8p83T9rXJWkz0E0rDdQ
lGtfPiB8HdgvZ9faG37SlzpYAur90Z9YLO8RBvFa89XJ/W1/CwFv03u3sgVDid1gg0brqrUkxPMt
LGVYcio7SMCDStJwktcsORpBYjyws79i1cPwKeRtyugUxODU2M6pgSXj0mwY2cWYr7zA+wCnjNfS
xZKQ/mtzJGMOz+UqDKOIlAj6zPc8CmP5a0EH1d31u4Js2u921xKp6RIZznM9KnFE77KT28vZxFFO
jeZoDsSimDO2dzlbWIQYuY4qBdacdtAHDJCmJmzuwkCGiDoijVrfDdoa3AQ2L080dklx5idw9EDO
s02LwIM0LPqSwuVJaqwCAkcM+IkphpM0iEsvtJpNL6c5FTVtBNfjrZ0U7QojhAcFQLIdp88dZ182
gl9B+ist+z5CJaWLZ0KKIL5azNSlo5MRyrpDLV8ZbpidpOu+gAP2SNt+IqZE+/dlJSAJQSUfz+iG
GS1XHr/EPVtni/bMAIHpIl3h7Nkx+nuglCtmhDstwJMQI1cwBZgTV82KUdSz3frorfsNlyz2E+K4
+ZnxeDjwZPRJQp+U+Ym95MspSToGgxVFX/ShlOKuzW1uutziQPSXf9pQi77Oe7muhq074uYU+yF8
d+HoOJfn6niNPKDeN+DzZLDt52FUashNavN75sv09uu1dEiYDlec/T1QxPa8U60f/jmj+65vodlD
k4EWtD37S7jjm5K22Mg8iCSpjNQpHBcJ6CjP2WBKWJ28JIZLTxfJMHVfajx7sMgTNIplIvMdqPFa
Ne7wLJTRiktaCMOGt5On7GavjVDbNkAT/lj+QSNqoW/ENU0rcVArDfb/0UvaOAAGFDAp7gelE4/l
Y5fAOLueLwA60SoVXSu2ZXNHAsVn3kuttS/Lu4pgEgD5wfLbHUtncmU/rhjBatsqsKIk4iNfAFis
yYmTCxxZqOYXEE1zW1ImDKdva80RkqVOzuPlAmVH5V7iUORcdhvMAtZ7mh7G0oZ9KDss4CG8WOAW
tQA5pl1zVj2i9sx3fA0/2emPyREYS/961BQE92i+GfzM169ybZrA1RoCXQEoyomsI2yAfX1x02+m
KezACPuHfVTWl++CQ9cADxRzqaTc6K4+AED3ARftctsWCSpgo3YtvOqeMMVrACw2bpKSofhT32fh
J84GjhvgI8p/WRtto63GaEif9sCt6Um1Vcq4o/vANl/s3GTWfvmtx4ygOWIr+CxFNtOu4LYBQY/+
FKyu8eQv4Rstvt4YV9Hj5HFE0uZK35LLoxuqKjRVMO/l+Wtcz6YxbrnITvwuIpodlABjpidQlEiP
k86/2hm5qG3HZxZ6nTjWeAjMs/2EHJ8Iz5eBZ0jASI2xvf8smDDaoY2HOkWb2LvGXGHqyQZD8Ard
ecp920dn8MX2x1RvRorz26DtFH56IKCFlXTiE2wo81lAUjz2+rPBMRwaoNC1BO3tzG2fjnrfbo09
6UR+QzndE84ck5efSDWr2YtvZZHu8BX7ntpHE6l4Knc7qvo7uHf9z0P/RngPKjKw3U0abuSkyafG
gRxyErhY5hhp0kBLmHdLyhFElhrlhunaHqC7uGHIQVO6/jf9KQtYcH6UxC3YIKKm3wGPoqVhEPG+
AwQlm2xwvyEuUJP6PdXLJDgCJoqKTNmkypDmY0Vy1EejIfjyjChmVouu3A95mVO8gX685iAcNjTI
7vIjPM1ky4KdgRh3GHyA6/fP6VPUVulVyX7RPUQ7RbxnEfpFZ9+dHrx7kFxBXUzapyHC5+aiLKn6
de3uKazlIJTpN4gfxNLKRGJjU4yyMfjaURIbnW5JkXBrCxXQNGvP3TvFDjVN51ISpOmlkYv8YkfM
aS7DDURdZVjJcVko5ATj49LCzpdTGGsjQuYVjl5aI5JNgVjcFRaTSUKyrte/2uAbzz3Tsvm+cwCY
ikDuqQX8/JHa2unzEOUB8+bltgF83pSl5KQzJrm99sRYFEwgqx2m8FDPdLgZaMswgkCedmE8hJua
pKG9cG/NvQU4lhT3VCIVzZXtu4KH9RlxIa3EJmBIgSCrPNLAVhsgv8Ui1KBluk5+vzuRTp9xQ9iN
JEKpSokOFx07S0qGhwz8Her0Mg/AfrDohcw7a+Yt/ncvJF2bhUxabom85pfnBDazbYVQlrbHcsYJ
BbvC9fzBRIjZG+kPuBxUFPngWT52UPO5u5O9+HgtEt7t+PXZMVwl2HzheJLBGzkChzzs0uAKnsaH
5bU9Z+zuK46vYIXaFcRdr+Eivu2PIBGiJTxkDCGnqCatqAxCOojSRJ5YnQlUq+dpnjjR5qp72Vl8
KyrqR75WO3UNAOLmhPqWAdVPwjW0s2SuAJLsbo28Mx7KeE2q/Q6bYFadFmtLuxXKqYjVZfCiMP5N
WlJARITsx3RjEl+FZiDhqGYvQLP/vP2fNoA4YcRSqIIPmmbmcoMGT0ZJ/UVoCdx6Hiu+AMdyuSaa
wUud6SgBSLkaOCb+VtjSNASyWuuFbYfNywpp7A5Cmg3Nq2YXDVjob2SSs9mgpuIvrgXRRCZiUlNN
z8Cfm+73Xt44eU7RPgRWbZouRpaqY5dohYMMlBjHA02HYsChYIA49R5pmzwvtftCO9mgm6nlBLwU
xGndmHqv+uhDORIz/vY0XPwy1R8C+Y/8rUSpouEZ3pG4tAZcwwuCz9qjR37kvoHvODeSIfvuXr48
qTyDkd2rV307weYOzYncwknMOwCBnqYpiuaWH5Nu+oIAINLeZ8+QuNsjppw0pQiJm18Ip8E6MPJp
LJHUizaS4JLVA+fsxdbp6raYb608OdIDf0j1Yr+MW7nVzoUTa9+ve2aE9jwA+x2rKUTkkP3FH3Nt
Q+/tIW/Y13EdM9SZEpio8mscko/Sgnthun6H9lSU66GkbIy6F660Pi/bB4YSUranlMzd4sBZ5DZd
143INc0byOxCZqp9kSGLtcJg2xZt/wwWwgiV110opMfQq/Qdl5goPbctu9I7l3gf6lZqgnIMoDtG
hsf2icR0IHzvHeMV8lG86+sCrnoFWu/SJR3suE6ygtzVQpdnExbn2C+4GGcT8+USAW25S9Anao0F
KDk0g5ApqlSrYgEcQRFOBfjWBBSulREppALPBv6zcbp2SSKfggvcKV4d4xlA07qKAR/XL8hcg7rK
iSx5gGG5EEkLow5/SAxv2WSmtknqTgUmxxR3G/96krtFdMF43F1ytRAavLoJGJJG8F/El0iUs6/D
g5fPiMPjkNIw+3htCN6rtMrbmtSa2fnD5uJuwkbGvH2oiTQlqigpZ1pim5R9czUhLJZKiaogxNXj
7cY+nk4U0RFWcMNYf+X9A/o/7Vyo2PUR3B6r4tX+zhOO1yHQCEy0TzZ2OV1tZxEOB4KwF658/faH
7xPyGGtPHkLUrpGrn7gZGc+mKeJgIodYTVszv2Ig5yISDmqpN8UgdxjHTzuyPjfiDUVrm+gZSsWw
9NYAWUlFCBcxrfaMzhGgoypbj+CQgH9xWD8uak+ZfxJ/yfbTLn6hYgyh/duAFBsrE8CFb+HwdesD
3wo76yvb8RP0isGsQ1k/zW0tVF8RWgKp+CA2gOyr2N+AnCa2O4R5wPR6emIVZXa15sDlkaLDwEMv
2vCjg4SnSkWrjf6gsUjrwWAzaxukTvyjW+NEIjzxbASKP0EpBG0EJMlZD4A6WH5Oa2i0Zpq+n+uh
u42guOfKmEKHzXeUClbP8tQ3CtnbiLwfn+vRLTMCqP5V3AHnlA9s7pPYxFxeoofKioHUXzi42tGq
2YLdsfJnmNL3mXy1MUsr/ejSU9mEKfiK4xqQEcvpNX2RsMlxKpKstOcCv6eMkr/Df+lu3WvV3BYa
44TJevYTxy0W2DF04cBJ9G9PjZNcNZPHyn8aeEpLjbVQy8z74ofLh8X0HO588K55yCedCZVumzFt
yvgf3wSPGJ9Bg38csATdK5Cs//iXBhKP9u2Yy/rtvCmXTKywyfSHBCe7cS47rKA1UE+zW+cV+kqn
sPC/91t5gLegJYe0FexrnW9Asf0jXpVzRFgxNhEwjfZiDrHy0qkjMOWDTpyjzaOEs1rnCUzHucDD
AKPC0dCIz9LufWAfjiTqUphIhCvP2JDZyEkLBuZDJLSnkg2W47xGoxM0CeoddxqwACI40b40/xlz
5c8Za58U9crvqum3Okyn3k8VHE40lUZoL2buFERvLZrevHod2quxuqHCt8+wMFkcf3W1GLIlxBcd
YJKgW/s5OPgYody2sDZYbKA5H98QrpPPxnZ5SiUnE0QkLlxCz8kKVCbhnG8RttK6Iq4KfvQi/9H3
TGY95SzfvILKvh6HR8Ye3XbLaa6PXVVWFGJCcXKUkK60a8L1OMs/z/P2lKkrbxF+uVNzHb7KS3W7
o0zq8v+7WUIxwWU5PS8+esNdyQLGZvSA0SogKrZgISOu5PSXkGZ5meg/04VPGZGx++GhRm+T+0RC
SFfiu8kMhbrfRkoOmgj5ssq7/W8n0iwp8mSkKzGDeZv4oZDVU+Tjn5WMtZM3uIXj9pZYGEI0ZAyy
9e/PCL3fcJ186d3mvpu6wNBy0tYKTUFk/8kOj8xqmdL291XCbHRy4jtQI5jRQMlafpmPPZdJErZA
U/yIO2CkBcc0AKnXsOdxHYQtGB597qsGlcb5lcifGJtO0tTv7CNxODaZO7+M4ffSsnkWXS+pstka
ksh+ZFkp3qlMRyNgwR2EGcHeu+KWT/cPg2oFxuKleiPJ9Q8BBdJF6fgeamcsVU6W8LPlJWwQM4BS
VdlYnXaKwtn9FjVdBoFrfNla4WdvR7xC+AxFbHsJvkBc/v6erIWi8nZeJupvsyKQ8mifnT1zU5L1
0fTuFaFeAmjeWgOUffdxgKYdW5Tq8a91t3rNCfoT5qjU6+w/DwPNxGuWYOZK4ZtSpZtYYE9o2TAB
nGWxTmgzJQN2H/6DZz7kNBE76ROyB/yrsexRNP7vI+4Lo00z9gDoojR9WXJIF5eNVbMdPl5z3c5i
2/xl/2NaJQjMRiIG6yp5xpFM+7e17qSsgu14C3/LwQKGyzDQfOxbsGpyJLNGdMBxfVDSGpIW8rvp
LCX2IrJdsopZxfj7/sx7FCv3fFIujvvHsCsJjDEnwUkhEuHT9MqEC3pZJaNPls5RKt6Vu0eHF6Br
4gSkAqvnAM/7apId+ilwzAHtjMGOovpTLMce6bfqXb9lbuptbdaDbxR78cN+SDRIte3JUzPzbYI8
VcfEhU+POqI6pVKJFIKEbtma9jGtCVT8wPljtcq6Gj/lGJ5r3iVDp42uT1w30B8QBttPwFz6n4J2
G/di/4HQfMg9TkLRq1S83RJ1+dyLHSQQpepKJ+OCwv5fkb3H3j3Y3PUAeZDLaqfTdyhA1lqBJjuG
g9sf6B135XjH6k6INDDmAd1ZwkrSKsWw04pq2QqXZG1s/9638VFgmUTG28E0paAZs/bnWlIz2X2j
LW72zLUjbwd6K3MOJIoqGau+tExu+ATStOkRuS9vz4lPU1w7YTaL9T5WaSE4+vQ2TpIqlxuiuFcU
SrAoXeRqFEI270ol0izCxBwD4tBZkeaLA2u9ScKit0UOpFbZio96caIFIqtcPRLIFgfBEVkb0fyq
n/3luOAmIMLfzRqE6SysV0Reht96CDQFkBewoMyYlTaP3Df29AitB69AC9VcutXZ3tDDv+2BakfS
rJxHrWY8UBXWl0Z4gFhSp2YWJBVsoYNOXAh/vUVwL2VXZVIQiQPYgimPCzLLaPa6wHgS5Srx0lQ2
mAfL2ywXoyVaeB7uZVvzLNwICYUjEpr6TF42LZM1J8t7nxyOroSPdDiHiscAnsFGm+XbeF2fgO4M
dFxscLhjcik/ev+75geZvwAvbyK4pjIHKFAuusN8RdeCrEDImL+7Z/GuGpnncQrNYR+02rAYzIAN
7XPmtIQdZMC4HOQcGGnstuuUgSwuxx+MWtRNWNCXuHH61SsjzBDHjsI1qTE3S/K/NStsQHXqTbuq
VihGOo2hZpK3khJtbSh/HRotHsRaiZnuJVyWmeCDfop4isa3rOh11qPKEEC+zoPAZE/Sj9+Nemsz
YwYKzL9PjCIwdqvuypE+ZfPSEfhmL8ULpphtBj77mzb+8XWCQeMWo8UQvHxoFBzuvgxDEl6LftuO
j/jIeDKtdsh8VTXNcj76L8YqfuC182rPNz0ejI1u99oFmniicYwOX7IqpYrrFurzaa0nwNyZT9BW
8EmUt+jkSwHN2VjMuZBnjUutZS7tM/3Q2PkmIJEVN312JlTw0VYiMHf8qUemMgwuilRPeeGoGflR
atzD10lMQI7jvFjnAKO7OaNyJiszZLYByh24dQVbdS/ckk/NDDS4WheqljvpdvPfzEV2LBAG+cbc
Kp4f14DozToPNGREo+x1bKSWh2ouwoXXZuH9lefV866XQp8gonztidg7UO+cw2ays7W2/Yeq8GDO
0KbHN75nhBuiAhLMVrIGu8sCQDn6QB/jBkIsjfvvxRY85wPoettei6Mh9Q9M7hMSfu/0nrCPEqPb
7b/BNcFwhfdHBcDBd8NkcA/BxOSUqOdLQbg65azStrrDPqC5yYnA/6XLEagGhSJ5tD80UFcGmWyc
h/KLNdEoYrSo1rQ13sev0h9/QJqpwvOPVSc2WhPfvrii9LOyBkGUiR4zT6321MA0/AFPo5s+hzMw
zO8CL7HOdgvkN3vOxplEfHlwyKpnxiIGCMEAH+7QBcSMKMmNMY1d2IScAfYtM7VoXn5iEEM+IsU4
azJgxeYcPpM5YKR4++9KrT0NzShS+qRobeS9/9CBtfvEjVQwP3hIdqgeOiGlE21irxLHMMagpYGs
Sffrauoe8USDqCqKO9wqA9bBcvoaO/qLNI11ROipx554Ivg6XkXf43dLsSdPzBrlvjHF62e9r3V5
/V9O14IEWtZJSWh/8xEbJoLQI+JEjgVtX1ONYNpRmpIyK2lw6FyHSS4/Kzj0FXyDcpn+jbP7Jg+5
/b0/TK9iO939aYW2XR/IKRm2BZvCWeLdFcmtnXXA8g8ojsZvEba5QvgAx9cYzdNOgAbdhY6QzEgE
//Jixte1t/V/oUBpT3AeI1w0CSYx+GrEgcDcg9gEN//ReWaGWYCxkCdEE/2NhZW0pBp16paHFSZS
IDp0xAgcZrowFQfi5O5d7btVCbBuJ8OwDgrDSbOvHfu13ejOiLvfNup5UKuz+k2jtZpLceWj8i7f
cvO0GtU+jIypepo8Wf/8NWKLFv5ev78RmrMcAvc3ns8jclK9j7C6RF9iDc3FMnN7PvVdMYT56hc7
wlWkYjy8wMuhhOO73qo/1fqghMhW2imRw2Mrd6jsQvH6cj9xarnZ+1V7v47eTSc++1xyaO1zJkEz
aJMu+Ik//pINrDzY6UJBTTn3gQMw0jyQRTZ9VOcg0gp+fsQkmUyVSwr6j5gO9Agw2FCEaZjP9V5i
VvtVokSK6S9fZpI8NoDDIMJ2Bs+S/s9w6H+MDjTG6V85Lv0nNhBOKU+sDbofNsKWZ5qYpqpE4JVv
Cz7BDZ5y87rVV1nTIUl0O0oSfyTG8PztaJo8U7q1/atciVCS/NUUc+ws1ApC34uLRsXviq+S5TL9
Qf2l4PUkqBjw0hn7hO1m9aX0l1SebL9vMDrcczXdpmGSb28UCQ3XU0pfTbGPtWdRtcx6LhQBHjf1
sxxyTmcueUf/C2nhcOiuW2valSCDbYOJ3RIfJjU3OkV3sUR9Wma5WAluEe56Ywxkzfr4/aVw9Jxy
mqgJqfgRhFcIk7a1L72J8XQ3+Qma2/GcCCapDFjVl4VPFn4xso+0hbhyvnK/iVktSGrob8VaCs5j
X7YtQOOCTDvG2gIBYTl7K7yEMojhFGq8yO+h9+PcA6GhYkRrB2hsLOZqlC5vcyYiHH97n09h026I
uBTv/39poGou3qOD2Nf8wSaSt9eLrc7d2RSsATa5pkeiA83aThL+fMjm0dgSSMdjZkFQLNOnFMVO
JTI+Pof2bGHcjiFK8PeCKPzwQY3mGVrHXsUMOrpfSaxICXWTeVSAWdrP41TxA/mFVLSi3aggnovL
gLC78Sp36ve9TYhjAUyPTbkFux++SkhUf70aZ17pbLTds+wFSt/OLRuXOBGoaJqHb5Htst6MVGTQ
yb1xrgakuT8Nup24jid9D2cYjqYIV63ivMHc6WklIMuWyUo3JSRDbz1K06YSxVM8mxeqcMGpd74w
xMVC/7fTboml1/Sb+lwe4z/NlBTjYc1nOPmokK8RIu2Ic5CDT9EtkJYh2ZvCGb/WZYPtlxsoa56h
6yBuRsdaPBzxlddLvBwT0YoRI6IAfIrrkuykPFcdb83Q3WfSdv7SFZvBI/ERAZ7PAVbY3YwhaA+h
VMpZUd0BH0L9ErqecQ6fMBQSMJLjgYYfRH5sfXrUdd+nxZ+O8nZP4wfjnYEKd/0mq/o6Xfpf1Spe
gJxflCzvQo6scNy2QOCLR7WwbvkDn+9FNduXKCs7sXpsgfH8HbktUZN0d9f21c52DjdRu23iuoG6
rDo/r0yqa7tfVmRld45n6Qip3OQugP5wad838V44oWmVDgV/nbnYTr6xmoDNS0XIPnU2UVdcvtOP
xZsB3TTY8KVi0wM3n4hmOapYxgTMg1rC2bLEyUfHWb+1KqcfXwv+ThDKdvBfBE2AdJBRlIDe4uLH
jkKuPg2XTcHrF8WlB7a5OSVx3hO8aKoNqfPgO1xSXBn2G7FPMjZyY1aAmzr7lTaffOARgXuX7ETi
0fHXo4Z0Z8KjvAW3y2ZFR6cHmIgcPHzYZvpec/DV4ee9rIIvI8pmkF5kF678kCykZ8h1Dq4Zfu1R
sFaJmM0s7UK/aCZPYfTUP/JVRTc19QNdctRkqn1MB38sq/rp6VDOA5di0oDB/Xm53HHKlyv6RVO2
emWSiFLALXDfUAFPCuLQMEcu6gmyPHyLK53WEELH+Ib58/hTAjxBVxtUIMOPJyQQV+Z7MHwpqNds
U9okqTKou8/NUFf5YL/6uAr4jdvUKt1BVdO3Ir2paPqZMLMhiR3YnhuHd3uTE2XMyOdNNQnDN0Uc
44mwJ2QyxiHBzepzjf7SiItRU7D5AK8aH0SFg/rtDeipr9Tvd2fw1lReFNDjo0lCpnU+VC2HRn8C
6IeP/C42uM1kwcDf3I7wo9zILRbTmVZZymRC9+yXAeMj1RF8pmlFWbMjgQ2Vn1eQgxrw1XJFgiOa
TwXzR4/M+Q8t7ccFk1Z+m98Ns9Td0ZURCRK0ifBGijhSCuIdc2TxK1zMLw1aJlS9dtHfrgqlWplZ
fkNlAkmEs5goY8yc5uxRrSFwZlPU6T1Ma1S/vf2ZO/Kt2v/qrYuqjn79aJN/JbZl+CThDEdc0w62
gUym3fYSM1gYbQQE8N8NO90rExQZuhy7qykzSRdG+lRjuv5if45h1Q5cowAeE2oaYwzmfRomTPd0
k8cBDg5AZ5trakG+AyjorwYsgxDQJkQUnmgRJ+CRn60UW83jT/d9Mh6H/vbTPkhulIToC7eff9tD
CnzCtH+vS1omNFlNl2vXsyi1h7SOj/GakWLLjfcYItIBmA5vVqwTAiQ+2tBP3qxtdWhDatv6OzIv
3fX/lTWBzVGnGkxWlpS3GLNLylOckyvOxAn0LTnIiyCcB4InxHox6xxkAF4DSEmg8E3w2j1AkR0O
iDuYTJBJ+Rccmlimyc3SMo/c2ZOrDmOFQQ/aG4yqT91ypSIf/+LTr8tNruCcRAjrrEhBKQwleTMu
W0BuORfeLNs2J0QY9IY0/Is6Kv5I21DuxGWmkIGe/3XpfMGxpRHYZCoXvYHVZmX3UopX4Rpbf1n3
RVeVUWiQKN3UxUE94rkoUqDt1YQan6p0Ih6dGwURPDCwGxofJVodYNBimy+UJ1G0j7pIMiZiqINc
ptvJvut6UldVKyDsnA+WePF1SHPziwrse7uh/Lh9t3hDCXYcyblf5/U+NwstSsJH8O6udaJ2Fuzc
7P0aGtdBlt7yECr8no1Wpou/dOwRTCWj8jnLiE4/QdiqYtj7BplONTc0O1qVFW74LocgfU6HPHMw
3djTGYoU/I9qmgd0xQu/3vxSlvnHWSdI2NckREZyZ2NsZwu7NCWXYSdOh2JMgMM0VaQvy11D9aWn
hEh52szGhjEKyeX99C+lCWsYWWQqwlt4m3EALjmnIR/viuIafevQBIRsMhYL1Ht9h5Fk2IMxo9uy
rlWzfsTo6YLl6SvWkP0NP9QOzSy2L9yZvs3BofJPWZfjGZAq/diWSZdhumuk06y8DND5le+jD7LF
YnMv8E5i8n7BCOlEdP6FwCQN9gVwu1oPmJ9pZ2ve7FOduss82z0u3/lea91dD0AzyfZcvE990SqC
FBRBilowMyj9+vYQmSpvZ1eQ79FO7HYAZiENAuc7TNWODzQbhdXf84hSREdl+EWg0W2NfMuS3wt4
KsPSatlm3gYFWt5h/EogQwY9CIov24ujHY7QsIGOsiLH+v6U+fu1sDHZWsNwKXgnf9q/TJaMO0Mh
8LG8mnccumz/3SK59LrRuDWPdk666PonUI08O8pWB/4dkpE3ixJ/2Z+pKeQb3j4/PVzWsKm1qQnx
UtjSRxX2eAGYdPFGQzO83rBsTcEo1VG5QNNGnpyUC2kiOGStnRRsHpEetagwYT5zAhcs2QwmF6OK
lv+NvObMl0mXMmEgx6xS+MTV7JggzNv5QA5n/7Z+KH3C96YqwM//gA/l0VEmEZBFDubVvvMM1j4W
TbNHgVGWUCbdcreYqyMHqZd2jYDdtS6f9EeCcoPppPiHQJNPSLVZnZpj9mm8g7uQcx0DbUu+2FEM
Heh4f26hIv6UijRUmA5GQBigXaSqwyGGVaZkpE+PhR9jRqDIkHdpMY+fy5GLjuuWJr9CVru2vd1f
gg5jwd5JA4sXHxcojZe+ilh0GUJxIjPl2xjwQ8LG6jT9iE/bXqrXxsNosB9daCQRvodtybHzeGXw
zNLU3krrBhzyKXmtoIRY47YXgaQzsQHjso+8FXVh52F+iNOHNJBgnmPhFcNL9hJiqn6IyEJ8kn8M
xlE0jrXXaaTw1Fg9DhMu7ROq3C/jkPHTe9OT9M3j8A6In8thsum0cSaWh5d9nwK7fnUBCDjx7TO8
xVLQyaBjL9PFl3QtDX0vsjbRTmJOgU6wLdTeIh3lUD5vl5QpSSREfoFxDgyqBfUpV93alacuwUGR
THmYMZOjohFurHag+2Zm4J80tReDmOKh0hwO1DIUUahtQl5KwWd21OIdDJJcx3bKQ5IM98w0bXSk
I27PMDFuLI21vHrCfAFGwofqfFCXkX1bHgzT+dg+C3DyxF1Y7+tT+SvaD4b44xcMmK1jzDhRVSIo
mX1NA4aTUvZKI4cfhfpkZTi2BENoLiRFgxx+sgoMRnfFOCyNIiGhpgZ+8ioT6a44SaMzDjPY4MNH
k6TOav3dR47dDtWm5Mc9bAvo5He59dCoz7/VgvzkuRii9ZgqfQDPAGim2lJANlifGJaXFtbomvHm
ywgYz04zp4/hIGjb57qHcQxKS+uhZwC6w1EH1Moq/FXMwzXmsoTNZfo2D4vMruM6YU+6LcJLmGmc
xjq5b7Dsu8abFVRRNiPZ9MtO7lwZOhkNf7AFV2iLh1W3F8szBNFyGErJnQTjqpAp14IFfL5CmR11
ow8a+FxvOUkbap3BdVgpIF1iOy/1Yd8bkGm9tyuF08vzeTNkHqfoKBP7eIIfru89t3jaD1cqHz67
s0kDZ4ZX3/Qd8/Oef8kOt1wTCqaE905XCTcbhCq5i9BHLKLpLmeMVBcuXlU7mSdpmkMjv1BnGQ8t
bx5p1wH7lnUTTTpL00dZn61NeEm9cMFQThXUrjXQGqbolSf+xdM1oz/Fu+XmCiVRW1O5a7B1lipw
vFAKaHASm7sES9Uwiu0mwzSDbvCFLHpiDZDY7euuanjVS3tuxRc0bkHrI/9j0iCR2PCgCKqCLpn8
7ZCNijvwAWQSoqT2els6+lxEg2OhP7lq6bWgdffNFb++RyLJox7Q7uKFpnbmlMiSanc4FgIOcPFo
5nVU5XtB1/Fo4I1RoysHQkFN1z/MgPZwAalLcuVqGEshNVdZw+of9zBfzr0hti3arGHeQC98xBpd
iXhtQtQMhskIvGtYZ/oPOC7a8rHmEjYOGgZRllCneZG2BaPPKMqTeoewjnbhElDJDiQEjrTJ+zIi
fr173YfOUIiXk5U5zjXnnDsxfVxPyeOZebsGPfgB6s1Jo6AvcGU9PRAj9ZxzuKo3wn+Rv6g3m8A1
844LxsAHNUKjLYdUpRa63oqna9j+kSa5xQVgOm53HGOlN+D8mTZU8te8yVRgYPNQLDIWazTiyE5h
73RMDweDPVF82Dzke+VG3EdXsY4ySR5X4n1k3cK2CRbTcVVNJw+Xkhd04WJPMxhm1Skaho9PGSqb
Br/odXPTseQnYoxj45gEamg1wuGzm9zA8YRX4B2/4bhl0P5Nmqf6jdz2M0XCFHIHKGrzYXmsyH80
vAnJhN+lRP9s2tSJ45427mZbruC1C8cp2w08uax966/EFz4VVkB2euWJLAv9eZ40Hqm4WZDwntbg
H8fge1nGVss4B6RJIkmUjIeiSmxEyDYbKqYMMN4Qf22KugSlPJkTi6Ok0i1cGVTw/TYbpdCKpGg6
hmR/0DNdsV57JYjnwz/MsHf4tUTgtvsjoAncFq7jOObMZh9JRh+960Jk5q+xG0fVDakb4Sd3oSeG
q8HDwfLuTRjpTtxId1PDlDOiwyEaOgnoNxhLYEcwaiP5N9UbyYiR/jbqKvq5/6MQF9yBZ9wSrIB3
0oIf36et7gijw4qX8Tsr5/NtFSAN+xg7WBfiwWtcvOBPiq9R8jk89l/Lv9LRNEWogHHu0fBAX7SX
PhZrTHdgArfLyODczeOh5uVtj4YHEDWPTyhNMcw5FF4YHB48bOIb1T1DofNS3hSBpomXrGujv4BR
wIxUuvNrIrD+kGeODYFYBeLg+MiNl7yVXhSsIM+eq/fnzI9Kgzex45KjIgyAKiOav885MqknKBt6
epm9MkuUmDSKrRBrb/Ekc2/Qw9UeOk+PpObE8v2UAY6qa+SdkWwO0/UOHptAOnkaRUC8h8DRd+Oz
egHhkAcPHDhOUKd9agZ+T/2Yh85ewxwQMOwuYB2gkO4Rx4NJM3zetremzgR3iocFo801sR5tnapi
Za7xgi4CiVudQYsFn7zby+TV6terNkiIr+gwMHQweP5AigwTl4otzMxk8JR/JGT14If0fVEqHDXX
t9Kk1NFpmB2e49iPOLEgt9VCMWmpE4J6D11exRX4kePJKJqhY+nH0x433p9toymLNJ9TpzJWdT3o
VEIwtO/CoKN5svRTCAYVcspfLlDaxrbUDETJ6zIEphxBJ2K1bfZceH58N21syqzn+gBLTFeeeQkz
NUqW/0s5WMGT7jK0YdK9Kv7GLVDRIbjlbMQ9pzr+aXfKxgAbfFr3wyPN7zot4a3gxR7AzfPGFhM1
fGQoBTPOKm9fLb7no3XW+x8bYm8u63ebW3nSTR1JfSLLdJMomF7t7BmzFggTpFVh1v53xU1f8qkX
/VoL6wiqdXf0VXNCiHcCbeQEBxatUwdOtDsk2fjGxUgdBrQQZA3rgZpNXWcjv4yudfNsR39esgi1
p+YxkwfOXaNsIkF29bxgKgpZtKsjfrR+80G2vJEKvFQNsdgNl6e4hX3TTyLkfJq1/srC/V93xBaA
ujB0KLxIL7bbJWLCy5riB62LdB/UGYAz/03+8XqdkUzVxLilI1XzdMnzzk5+0RdTS2AxbQuhiQ2M
MLOi/lZZYxPeCa/xQgE1Z9/1soIdnNbbAYuyp4uyNZ/G4n8808kJFiFZdp7DHeWWMKDNqM6vZ7Ns
VuQb4p4vicJku6udrJQbeSg/AIvGcWt5apkkA1MbVDbQqHPzKXvJjq61brHn6OS2ljldxF5hiFQM
KCFJgzYbyH43GKsdQGn0QqJ9X3HiMNSEjDu3j2jovGF/GzRRyhECSqY3rysMRbvcVvEY/vaWws0U
SdU9weaOcNuGHyJZm8JT4oUv5/a1sP8KPxH7e9vvor1eZK+txK68ydsnUn7OGvAMBYhs22eV5nUU
LLsaXAWUopvN0g/sE3eb5kYH/CjL4iQ3yz+EV3gHif9neaCVfvlJ/0tygfPnl41V16FuTvM7hcB5
d2pAD6bJpy+/HLx4TSwsDQABJ9cC4MOToA3HCo1BKfrGfWacJMErTUOoNE2qU7pMf6vZBUi/gOuy
WvlZX3UdFDdDfh392TGGQFAS3OkZUIgnFF2L9P6IxCmu2ghPj3zThJucbvu23WiUHiTFdpRkxw7X
L+kphuOIjL/6JwPysZsfvrZz26Vk1PsBaIr7SD2MFz0MaHcZYC0blmrtcIB/Ot5wV1Tu8Nkb4NxU
VhdBqOHEsYJiTzzpmdkhbqNoIjo0/O1jD8kgyQUHleXJIOI1HwkHlI/2cIFib60kmlr8AEaGuPrg
B3IBDBKda/alBewozdP0pAKDmJpMTkH+jwL60leIzBVYZ9aNxrH0nxQYdDJrTz6ktB6GpmWHEoHa
3mJ2wdr9I5gr4tMc++7qGFDWJphuzl4hwwoUzKN9EDlMYa5N4Aael8hKLt+lLW+ydr86kD8zw8hd
xOwB+lxu20S1U2hlX+bXQkFuigEAOM4fCkNSvZ9YYPbsE4piE3DHodBOTVUtbQ9PxgObdOeOFe0k
bq0Cx6bnLaArmIPms2f3FIiT2H0WG5g8k2kcS5I0/a4E5iqwnYTiX5RPChaPRrDqVraT4JkW90ie
yxm5OmfHnm8ntQ24Riyuhox4cOZLLsXTVUzNZdiLMcNvujtO5YYO0P3nHHdAhKIiijONunpN//7y
nLpkZFXw9yRU+dcYNQe5YFDo3wRfgt/7fendExbcugYJ1NVP1+0fCj6Inml0TRg2Ogpn+Yb7pyzM
0eds/ZYaRRs9Ev9zWZVZNsYsI5UeS6JLVG0leugRLrHoCgQBNL5u6m2A5Yuva3Ytmmf2zlnexKx0
3I032/MvkkTnrpEoTlRnBYak2b2x0ENnkSMM/gi1YxvWeI9TUTi0cruZy0SjQOfjeARqbauTvz7+
FfNNSOn2o4hBaE3tQ2SKo5xfmPatfT5eLsQHa22gF+07+tLnhMlS4hBYUqQJPSsfS/Xd1cY44I1B
3Uu8ouNgi+9n/ClgdsQ42erLJf+SGgWbBneYs6uGDMS3FkkduXYR/IWIrU5AOH69e21gmLt3t9bF
PUF88xMFvMs/ezuxmswFwbDCdnHxYi9Bha37qhT7FaOh2CHjm1HvV/D5If17uF3CdXXWFxJe13Hj
UiZCE7nWfP1/cDD5+c0uD26/1azuPraJ4UqxbmZxTnwNniwHHj9bXwOpIb6VS6C/+PjEvlEXnoQG
oR9bcJhPW/U3vec6Ac3agPLdzCP1tE8j3MEozXq8cJ7KUei3lIJX5FPfQ4/WNOikZj1dSv2P3Y9N
BwmzlvP8wABc+6p76ygCWdChVKZM1ezF8hpMmy9oQfY8S0xvz3NPWsjNdbU6dnFklh8nFTZgr6dg
VPw4vPTvjPVCrO3RvV+JkFLsHHbAD2OlA9/pAIst0d8E5U2FjUCTn1qjZIv0j5gRMXoJGuDAW6xL
bFUvpoUBnJ1sN6A/JO2HZSSXAB2gVbvag6dolZbUw+FbzPPUYx31fqPTM+asmzP/+i6lowqWEVgb
+5on0idjlIFugZ8Kfy7LBoE0ZECTkopl5kr1ibu/hapGrcv2Hq4e+PkYTT84+annduLYohIrEzid
LgulZ0ExCmE+hULz8sTrHKQyEFclvBLbqbC9TPzO2s65Gmd/TidMKRtQyZjttQL4fxGeFWqx1nt5
uPWFqy3iwJFKe+hFdO7T0V5GITQQCj5hHYh2PePnAUgK2fIv3jHksQKQs40/leOuvwOfgT0o6bcj
6EPPRIXFUaqhiGAx/yOR42q0ylihMjxxPM7ie6YTjmQc2SirkxFc8HU0jgbpATFXHJhYRvcGQEz3
lF6W6gwOhwuzNnR/l7imSF15L0TOCszTz4Z6gSJh/kq/N8Usn1g7P2pvPQqj2U+u5vjmXUbFX9lg
Khypd1BeX7ZSgyTX1+tR6dVmjXQUgSIijSizrR+5/iiEvx4RewRtnrEedqBxdVGn8I0alQdkJiHP
J69pa8Zd48S/SD4r7CZCi9tpnxPVU1fyXjz0jPb1LudfRD8YF+lNEZwDpzQxIz6NMpJEX2qzXKgo
JRELMkFwS6eLEvcg4U9T2sf+XQvbrUotUMIAfa9kHim+UdYxiuza6pNa7zb+kYVbIbHGL/K229PS
dXVHdAiMjkUiKSwvVQZYW9toKBZW5zV5OXh/yWpswppHNNBGY9eg1/kqo/bIqvC056CKUslKcqhn
Bnpn9RrQUpNYO+xG46Sj7vyh6wQf0RbRG8jAmRqdSbgIXxDAtESwvLzlHeMfOAk901QsYdpe81lc
8a5mty3B9Cwbbe82iuIi9dRWaI3sFwhAmlY5OEH+vQVfjFv9vz4WahUf8pQR0GHBHctzn5qk1NNk
4sdjvRt0N1OUqHRI5w+kMm3AaNy5FqaEZrtozlabUz7sSKSZWPl1KscKhLwhQfL3ezLle+wZNvvG
y0Llv7T/XgmnRU7W5q3paXz/C+9jgAFekYcWTJmJm3bUuwY7llvzqvB7nBONqB6nXs3VPIwvBZN5
cu0wbJnByrMx4ExKL+OwD0d1nYfL7XCwXHzUvCdKM/FXPb7IiANvCbvVFWdSXrLZSJ3twciP2h3m
nDQ3HthRtrZ5Cx9c+MH+L1A6TSBkb2Y0oTpRwc+mzT5sdA8HAQmrJY/as5xwbLGie9vKGwPJIMl4
5CNEwt5QmQ0mqcJPWqL+RRdgBOVSZkk3Qcx3BNBQpPu/8KP8W5XJW0nea3OOec4EIRcJ2vCVXXXJ
BUwuNmAvAzMXqrkd6vVFIv9BQ6hoNVaZJixBk7JH14zunYz+r8sgt5KZKKreuLMGmIhKCWES3FYm
YlHieBFAm92EqfKsO1my2nM3NXrOLZmWFwNswbrlmEguDv9RUahijfJhGUZWzDWbI3UJLQWKStV8
KL0z0zZc156cvuxUqU5p7ZOUTsexzy9bdp2hVaOt0pcj9wr2D3xrWbktZkmQihTm8bY8S65w7k6o
rYTDnQEM72zhKuBZd4cmCzTinUNT1ohgXd+vFpfMSMHlygS1Hjlm4eDRzdKQhWwBs+8pnNtHsq+Y
1kQbaJzJCmoZM657MjuXKB3HFcEfeGSRTe5sAds46qprAb1cMt5Jh2Te7/KgDvBoj7EYaqtPFrlH
heopa38k5X7xvH6beh6snI+B97yd0VuRk9RMiBizeje975TsUiNVRprTkQErIP2g+PCjhVSNJSt/
c5FmRdRG0om1GjQjf8mH7ONAMpN6ikbutUui4mEtYkcqAOJgpvZTmFfMHG3971a+sQUaP2H5sDku
HtntAMr6VPAApxJSh/rkLYmBLlOImt0j2+3eXZqoVQM/O9xBpqrj9NCtb/tGbGPhbVB9K5hhD8oL
7XktXk9LD/v0XiFGrLyXOU7/DkRRRtUuqiHwfwJHmeuil93lTbN/BrqscTkb2hvepMUR19MjvE1Q
lAbyCCbiOnAOa6hcU1SOH++76JDRnOV6/BOfyOYaRx+x3Nu4BovBghm2D2lNud5VOScoWeu2A6xp
GakIojx0S0xDZq992Ot6DO2lswL5u84l2BydQL/OHN2bDD6+JKfbHmAvaOJM0YiPRQxWaK5WLgSL
DoMw49QHFWzMDpiv6EX+j8K3B/SSHGh4LLB8r1uehHdCGEvR0M5MxcylZgT+4U2jThfNdTsjOd7V
03+3Qr9vl1KT21i0dbx7ue+xRkCiipJPdI3AVTf4piTZdHTXdc3QWXGsJzrrn7Yi/Jp2ki5Xs1S1
+MOnWp4VE7tFTjtO+GVgkvLibpcuBpjvS2D+76jX+pEtd7u0WxVoT105Vi3bxKfxDXHvZyGZbks5
LIfpYO96hw1X3v748p2I9ByYYDTYTFIlIRXeJSs+z4npmdYw0xd6W57fYzY7sdxmBnSqLLUxov6X
NbDmrD8PJkmSEmwHV/q7QhMGzpSwZtmO5+/Yf17yfHPwmbWNm1Xgx1cIL8dd/FYUTGC3vUdFBn6q
RtC2e7wuktDDNrP/xmFdZD6CmAtq8wRGQKd1Mvbt2mHJLXclnhC45UyxXHQKjbSaNwf1233YFFar
L2Nk1m4XpGNSQdWhntHFDxzSHEDxFhQs4itd40qPe8cTbeRNbTfpPlQKeNIBQAqQT020Kf/XnCvD
FmryyUDi89y5u9K1z74oZjxnmwms+UNO97ADo4pfbyt/LugWy9I+bvyyOnirflB0kuaoM4d3ed/m
PJVM10ZKBsqkCzE4IWeOq6zG87PtVFRlmy2BaUnKrMQH0sczln2cQXwIJtCJj0XavCBVMrbiKRM9
qALbTra1JRFyOjr3DxuH5vq6RjiZlj/4ybw0ASXvy9WiLG4YClyJuP0NZ8K01ADFYuNceVOY5FFm
wuE7KsS2V/rlv0AP832dactv3NHX6Kf0fOiCgIxxTICIiq4AH5DWPCTYEgZobtTIRfORJcLmTQrc
0tr+wd88N76FK+fc4pFEyTmXKc92Kl4P6+Mw3JMP5R58Xjp0/iXV6PkKQ/YyhXhqVwE8uak0Q0zj
RKVv5EMoDUw4DaHVkd3Sv2QeHC4uXjnFHv2aCkMbXil7drFBvhHGo8KC8aSMMywXxQHztr2GG9cO
4wXlWbXBA04Q+AoCEpvs0q9OChPEZRuk4YaUydjV6EkV7Qwd+o1jhFTz5V93ZT54yr/VgEs1GRYG
nBjcIR/nNyEYHvvi07d2NI6tNQihz8XqAkOWjNjhlPtpYYt+JpCdXSlM7RSuL3pHvq10doFL5RFq
MUHZlSM0MOCrOwUvFc8wUatDCYXW6ohcntAf57DOP1JjnjYaDmoSOWmKW3Tx5CVGUaVEAwyc97tV
PglWeZ0FpWd91QQsoRIuTFAvGB6/UJc6GgSXrVbVJgvVdxjTObnjxx7wGfvQ25LtlU1a9Vfa1hG1
XhHQmEq51HcUKPaSG0n9X1aG9iCjA9fLIDzFWP90YUV1/PQTKCVyFKO/kJIcI1/6F6splaMY2CNL
EUJy/VIhk1v85+yzSceiEiQZd042V7FiBHHOVpO/QQEhtoYBslf4D4nfGJudJxpF2l3cKtea2f2V
ZYj9ZgwPmf7w0Yyu9dbHML0PbZ4ucViMp+WMjSvxJeN/rvXa1F0Jof1NhgnF4yq2G9nbhTxjO/VK
SwrElRFVOQ0eSDVtKHT5petccgNKr0l5OqZ3e7OyBHLGIl7vz05lU1b7huLgniJhMps00wPeht0R
/6a1U9HecHtw1lxl2GtUQf+D+NfGo86rEbXPdPD7g7dT6OU2+CyXbpIYbqjLnuhdjmp2iuFrXyZt
+ZGSvo4UwiH1AWiFxfvN6bU3kU512/ynIWmLLvqhxiE2fTcbEtcRB2nlHC4I+cYOS/YFeMQPnyvh
vWPZvvFTbBAAYmmRIkHt69DcvCYMc77T61gbC1+7Ol9jcEceSoNHfJ6SKqf2mX7kho4Dfg2IyhwK
j/iBpWbCnUk3DpXfbL64lNgT/fLl8a4E+LTyS73VgFDQvSkqUd7/TLMgBje1KDYik1pOtOJOVY/A
ozrcdh8xkueqAeIMe60y/1jrdTm6Hgfm13spcjLcTRzfCz9ZWs52S+Lm/ShRcJAguwro17PS2Ut/
jmmMOpJDXL00xO/rzBGOil/U2aFYsqkA01I/PzuJwzV+y7ndpRL+pyVnxYBKib72QeTfJ6NoF3Hv
PGvaSHId4GITQEuQj2S6eyV6BwHbFUhhkrqvNggPOFeWxXmLw2AJSEYO3IB4mmBoqPcCa/qUaH1K
t/P4Os6RwRrS7ZkWn3oRZU9smjxqX1bniDTnF3LUmYPaRGvUS+g6WaljT5roIcr9jlTRvesRUTB0
C+bKb5OY+R5rKdVeEnqnRyWbIJtjL1JsaVcHJky3MyHPHAuR9zHG+hMsz9q4CgiFCj4fQQcVQDq8
yYd3xspVhWLhXL5FIIQATlMvHZ8ywYhDYi14IS9ltF8SMhiI2QxEOvQTsV9q1MW4wgkC8VzqXk/z
MMVE5yYdpA9LevcpcMEk8pVKZh7PWlNtLCVueTBQRvDrhBSQztZnYML0vjKgoscGfQUa5qzb+uQj
c7m3TjMtvaBbLqYX3cwSudaqgcgfIDbK3q/luxfSv5B/yWfl6GevqCd+XZ0tgY3g8zmFrcRlSPUK
lrx88gLXWH36/u15Btm7nmrSwZr+wI6+ta75imcynzPLaPk6rV+0QliWQ5gsVR3upgbM75D6QFxu
b85jflBnQ+gXD3G6bRHLTQxiYJc2OzSptHS+WV2/CNR8aDQS1cbf+aSpyv4o/sCSapCJm767ND/6
krRpxe7uiDgiqaZ1NQyl/fksM6AQZFri6uvLPJaI340eMI9wpNsc23Lzpxg/04S6CY2rdhzP99Vs
X8H8z2CFn3R8oKYCUhWnDbbQUudMxI/01iyu36Dm5peTTyCn/eV/CAgXPAafBcb52FIOgkpUUD82
9eUHN1dVxcKoA+AK7R8F70mWRxo5YSQc3xrEBMDNJFz9fuBpB+xpYzVUFj/DDbRGq/Mh0nXbcqxl
kToOLmG5il4IoQ/wt7ORpGXMg+WqYP0ofk+RLNHpzZV3Qu2Rzhw2BgVQpNuejNCMyX8wLZtuKCKR
FBd5mfQCUK1j+odjQEi/9YxM5cvoU6iYl/l4O+aWMHb3bn1x3RUNlny76mIzof8h5mWI/r0KC4UX
4FDVSu3FWe77SEwnQSU5/QVM6j1OnSvmhh7b3FI6EOHI7Gg+NVBKPrDNcwXjvBOXQwDxjEcr+Kzu
pmPfPo8BANxVdYhg+b4bRWHNJtkXpqaV+HY3x8Ps4e24xtN6xXhjGnW4mYqQ+y8Sa3PdS0pkHfkm
Q3emtoJxOrHYVzsLyV4+QPLftnomz7ONFsu86AKj05SZE8F4hx3UZnuP2yfz/2LOesNy4SCdfuXa
loa9YedvzwUVfNBh//16jWdFH7WDaobMGxSgTfMJ7L29asV+XE1uyNANa8VnDjupOECQlfIgsYhv
gOt5S7FiI19x+sycAPElAt0MnZOm1BkxepVcVt65RX47lwmWVonMNMePeCyysVv9+262BwaTMk+b
3LrRcVsrtp33YO3UkwFfopjd+1kydVsTg0ZqSUcJQi3NKMvEOFpP6KlZloEz7wvWOxWGIMWBXiMW
pcHn9hy+SYvVUMmjaHzqO08d+WjpZtbtKMoVClojEev+heWp+tAjkQy5e80/dbjVntaubIhsUzTJ
ZXUgat5fbkSYLCevfh1t9iRyOPSH3BI5RRBQWzv3M+DdqyE05oSZBfXZxpl0uidIBWkTZF+2TI0I
XAH79g2RY4wnNwN8Z2/ectcTdFqecWSBkwh0TwrfAbujpYKs0khbZ35eXfkcRBHnXP2ud7+Xculz
3OSfZoswhS3YQAd9VLM3FlVkKtV1v6s3+HGEcXQjOLh4yJLwJqrP6nDcaB9vqV7GJFMcO8FpYrXZ
/HSzuZv8pYyybIDFl24upwDzpl6D0FGZfQflecQVczVLOO+cqFbwOxRVImznMT5E/T7jllIQviLY
UMVIwRPu5M7wqIW6IpVIzm2AYSPOeLdEIeQn7p0MSNSOpzKZgh/TabXx+r5nfQyUf7Z0fp+ZmI55
E+fbF1WRvNaFy0MS5Dwy2hCba2DtoIfxVKL/DLTI16rNmsV4Jo+I9N++TNHX4n29SR7Fc3VjLH/V
3Jw9Kb2RkoK8dNzNHWVVCQNJrEyaqxDPomG6HHlip31QpnnRHwKnNs/GC1lk3U/DiDqtTWteJGuF
dtD4Sox4RWPSGvUbUU40eVFbqKl34pwqanxnxP1QQMRSM2B9Us0hgI+ks7nki0+aZUSGkmw0LqGy
DiU4sxK6nPs1Gtv5hag5YHoFgUKtX9TsBfU3NErYUSJ1tbzE3chNY3bBCY9lrGb1ud9FvX2l6Ttk
Mg/ErqxepaZxkztwaewiDcBzY7cICRxjwG6GIf6FG2w74PnMLcTWH9/SUFeab5jvrLfUZegpD/H8
svE0WHX3HVyvPtRsTNIiSfCeWGPWfAFlAHV0fEPshP5jxWyClKJ7tDq9FhdiQIqRE8usGx1+3xIS
WXV4TTSde9XD6B4J/xzg0UW2Ksizj95B8TLCln8/n9dLx4oOSMJyeJU5qH7VQ7UT7KZJ4YOEAMlU
kC1DXzA0R8jdD7xldcJwaS2eB5j1WpWZ4V1uFo56XI2ZfzgtMMIiy9mef9XCsTuZf2GW71jrS+xf
ta/FjBurVzDn8uCeaKGyGYJmLpwfjT1WnrGXITXeKY79px580O7w5morsIj4DwZQuloAVCNbseiV
GLFm3LUsCuGv1ACAhQluTXTzsdhmJJ+MSN02JfsBAC7miS2dRWGohYGxmg3K/kobUlsEUAQDFyD8
vGn5uTTJ+8EvGCtUchXQ5jEokdAK2PSJtGS0mQuSjPBZdgBlG9imavYqOr+BXH2HXOdfuCpQ5IA/
z/BOOsAPzrb5Q2ZUGWzZXbWnasJhHYvEfZiPhlh1fV6gB3RtJfiSSScYn1OrIpvja8n8bURmDi1G
lrW2dVNUWBFW6YpaV0IwnFhx6MH1Kyolt9ROZLJXNNyIxTtEGyQQxgFZOsr0lzESje+x/ZkePYFG
/2M3Ej6cWfUeYBVQsLCTHJhESW4QLQw9jgUrr9GmnkXNW5rJHhrK8xJGBFgbnp3g60Dxtc9cRxDJ
FeZ80Nr5BwQ/i3zTuG2Brx0DD1pXFDbwn1sSZAhfypu/ZJ8jIUxatheDruEvb/MeXNegy4bkaGdG
l+lrABbICunjqkxl2PvBn6E8BDmJ8a5fSL0PTprK+lmEhTBov/NGsn2Wp+0oLS52SPNPKSKIlZjC
rrElTgGN0dLNOtAJnq7bTngffrd2IcWPD8UsDzCfnuZ2tsjOJpkHiQYOp3XhT6SJUSQA8dCyoYac
crs0iOzKeMlVs1pq3Nt08topSUSoFsD1t7/fz5WtSF6OTh5YFzWjzHGmsAWVR+iJI3SYTyfatFoj
61/asKjLksSNb2HEbPjIJyPSRdeq8S6jA3vE+hxIfJfTu0EU29VD8w0gJTqW3Ca0PWbcEJkQaHNU
YiDRSQuRP661eouYmhu02VA2eXLIMqui0mMSFrEsygB6/s5RmTJLXaDAsQL3mznNqAgXE46qful0
Qfxr8KJJKSDZDP3/Pl1pYn+xPpKt8XEWoQTx6dWiVFn4q2mXQCvEHVt8WxKmg4XSB7pukYX7fYeV
zQ3LaUPLMQruiYYENZvIoBfEzaEoFQvlCyhPP6RTnm5iEeumqXjjOuOmBz0XJILnI1TFeQj5PpiB
ZC857jXm0WkgxSGxBIWnvw+f6uL2+A/vQTN3rJKR1wj1UQPR2WiMFVOmeRILXOmxd9oJ5ktPBT+n
DR3FrUHboYlr/Dij8hrozk5CspFb3D9Sp9Rwp5JfmA26aqh12xjpWu10cpTdaGPHWmtX3sH3Zh2n
3+5AwD5yghGwCRgm5FFBBOCprW9jpXTTzJ9wvDb80eFJKJMWU5w1+uFM/d2zuZw8MZTbcs+iRH7F
pkIvkF9fFI6l9MncmgdtoRSfuIyDGlMsQ+DPDBu02ziUgCvKutsqzKeS05PfUxxq4wppU3dnfdlO
8u2EGImBcvaGxHaPsz+0q/7rSLX1XoQMCzsirzg4mh7pkNLqeOsQE8EIdpVUBrQs39/Fpo+qz7Qw
+IMjO2h570/Sey+jEOYELNe0x48+idgWkLbZt0otYrjGz/IYg0RJttTheScpsQzAiSzJ92jlNZNX
9Q99zriCKd7MacatS/RTTxG4cO1dSPszmDjl+22YoEiMkaJcvtxpqOHvKhou0X1Kz7jYsbJNcN1M
g3ec0rpZNATF+S+pctj8WqB5rpAyCmmljcjhdSIIT7s60TYo7tqRrLmdqlc3frnwZO8Z/XSGMt0x
7I5FPjsp3MmkJwCg+W4jzv2MSL9S0OpT4ItmcBUlFqjFmCRZ4Zqeq5hp292Rawsv5oEDdNz2FbH/
SeT4Yz9Zi1xxUJdtajyRb542IE4M+WoquyFWXffzuwyLOwIk4dVNMadBHGkY7t3N3rYqpuPzxFTE
aUJs9UFreWBBf7nWqMXis/v0X44VYHrj7KkgpSDP+gFnMyiRVHfB8QQGriapmlxxh0ieyNNrFuEL
1u6upd92wMC5k1zbBaaeiMibqEdE8iVUQHruJdnz3iiMzImzgRxDl3IdPJdiX9AYTAdort97Tao3
l/OX3D8RtaXnUcHV7Ti27LM0HABHFktn2h7Uoz2mUOvMtdigIpddMBk5dNwiyydGpdvk0B54ba9G
4BXSTeSUY75CfGENr3uZsMLL7DGbMb++CiSzH6r74wlO2ZuTWZ/cbneKvcnsI32pPCHxcfGcjedz
PXF3zdfYw04Hfij2v4LpSvf0ST5oE5w1cx02boJCQOdAzBZ5+suzQBuXQ7iX8UC7t8XrB21mWo4f
WuTINEXV0PxsPo6a8/QN6z//v34BgOPlWhIVRskDx9WFYq4fBbiiaqm9NQ4RWIha8XPfzK5WAL2C
Zra8yUNY1wksZa9QsLTeyJnGN+FzJ+Oudumk08v0Fe80NBaO7M2pVbpNQP3P9nU4EXZ4I0Yz+2sA
NEDSnYZmyiG7y6jBBiFONTgfTc+WKrc5/7zXYHmoKFl+qvoqeOImaQ6yUqkCKcx90uNQyDPSicCy
0mF/YScJBcT69iJiMf4CQXE6HtmTVVppXWtJiuKygap/cjTgMH+b9S14GJQVw22MvjvcCCaQBS65
cs442JTCUJg67St5a55mC0DvwZHsPdbaIo3RJ2a2suU7NEZnSGrIiDKN1FqDRMhJk/MS0e3IwvmT
0ZCb0tUJewSaX/7NNbxyP9UBcBLBI7z098mFUpfT5XEoi2p7OGR4PKRSg3Trv49jg2YI1DApE3jF
njzUdbMK8itBLB8mkICH9XnZTjBniNzqp3J+JDD9oAfhJUmIsI4U4uObs5o7USFeanFEjZTGrB51
c+qjxcs26HJkCIL+PZd9b56A1w3EtXEVSRCdAZAm6UioWbgahjgNo6jFRvADXR7Yzzp0V9X74y/j
oSsUMXjI0LIQ88rIL4BzEqIGQlDp+RZp120oXdfmzYlwvvndsByhdS+2vtv78b5OCnfIqVYPSCzP
uBb4OScpYVHVo5NrEtbOX1ioh+aR29T86lS6JkUkY4DZ5VPYPxuvHxvdbExxIIIBRrS62aUYTnYz
nBOcDMffU5QhflO4cHynLR+W4iKc2picDeFKk3Fa70bQNWdPQCri19ocTimu8noxFk9kqrXtkjnx
J/eZ2KrW2+Tmkuzbox973Eh2OfzK3RBC1EU7e1TwmjxFERjz3ZInr+xaLdKEyrRDnk+zvQPjuDtl
QilyEc8Yx+thYpGbwgUikOU/Pu1F8JCRRSvRxD3D1Yn8Hcx1rVSyAMlmOCWBppB+Dex7kopVCSY4
9pzA4HG+gfYI+VxllcJ7xHgTYKlDE9p5CfBj0//yEh6PZzJxIauPy0AgTDJhGaFZ0GsXGy4lnDZY
KIsk59a9ddtsuEK6X62DtK1ZCgeqL4gvHrqPhxvDAQeC/WVC8w7mdCJca3BFjGQ1RN5atsZONKFj
zJ7DFaeCl5ncaxS2fbakEuxfBeSsVVayZ8mw1gOmFP/s+CTC0iEZqsPKSdF0YV4wP7Yb9IPjr03F
AerNJuyVIAGzaaJm5PUxPfGSfUptL+WeGp4/OCZANDNFIVbrIuYdCkotzfI8FUD1IAnmIcZnCixb
R2Gjno1YIL1SBwIepDVbvtv49Y/SNsWnBrMmJUXNThKe81y6UPLdm6dXme+jUFEDIYIkyjeTGY8w
LDm3rXanN3UgSPEOzKqQhkT4Vwn6h12e7w0zphF93+ro4UrgsLJpIru48LziGkNGaHFul2JuGvrh
xsEmH8WtBRo9e6V2gOuj77CDsfe/mmEAcJpeBP9Bna7lfudySqT3BuELF3FsDw+yB+xWm55QnSs4
ynZTog8NmKh7lMvjSUd0JB1ce6sr1ax8qTh4aHPrByiCQw/EpWTWh71f/FdOPzmkszabu6Qrw5DS
c/8u7isnpvxZ6ZC3KFk8C0jzaFEGS90T5SMTb1YRqJ7SS2TF2iWpPuMVpSbIyGjifNZ5sPL+kY6D
NwcnGu3blR73qP5w148/2DhRoO74G6D7+AJVounKyVVD5FFwesX39aU1IpZcIRQA1EtgBCt5+/O1
q8DjSgRJ8DofNMQk78BXtmNVerhCmh5fp//fEA/50oR1LVhOMYJw5nt4Tw2dM8rBh+n04TPq+zC4
0U0urWSEsV3GQFF5e5uEl41FbFYlBsY1KAok0q9k+2VDGBFb+aEdF1/v3tqUfq3tDrqncx/47dox
pg2u25olvXAhl1tNnDOCHK8wbaPrMW5MWOjC63AoBgm17uwOPYETcKXUJAp1DnW62DaSV8npMWmA
Tm2IBBnuB9q/UtF6eRxwg+rWCT50V5qZvJLGZQwD9s+tjVgUoDmJrmswj3nUGevdSkP2MI2gySgL
Xdnim9VWxAhScuXF+72c6ztYDOzjVJncoBuQ4/yIVlEYTlt0Mw8ygvAcgnki7fxU/P9S783sscbX
ewcaauyt/4OIFQVJtfYpxJyQH3AJLC+i7jEQiU/GjxFIwAAWEHWZMtA0FOfKkq6QWQicaHsouNVp
tFtzNuGaYJpEBxGfJwevyo7t2trk1nIN2KR1PPXB4+bCMX9OhJIy1oBFGC4iFmnnwBBGDzf5+drM
RFbMDLFLTQeuogyJ5owF7ufsKW0XUiy6tmjEBQh0HT4P845E70fpjc1iiFDC74ZDD4lAP/iOr6UJ
lbakHls/ZakAYXSymeQEWfHonUUhuMU8VyiHSOV/p4wwvleU1PHnn25yx4Qy79soVBFSP/+ceUZC
GC0L4osRr27+/sGos6AvrKjrEIEkylrpWIj5wdAADeS/eyWfXjFcXL/kQLgO5zEzr34o2HSKzfdb
80mbHuZ5lrdoqW56l8/JeviLTjVLy2Lx+8FeLECKJDq9TtJtv7xkHKLkj+XvMHW3+oV9vccxU0Za
eDvuNY1avGwdmzjQKIICrq7WveIA2kNEumePTymfWcdJvg52v1tG6u/66/DyaU2Cnd6lpWeuqETU
9QF5aHG5Ca5Lmd0so6jiC/5ueBNwG5QiywapY95QFpq+Eie8nMxrIBuGgz2E8ZeeIf9UWEVIETVB
0ZUnmLHwDQ87TgutnBO74i6k/yQpEKU//zoiaryp66jzxIiraPc4CWNtkOtCw91MMkxKsrPEGBjr
+nq8mZQjHUuVyCdnxGZJ8LwtL0rNwbg53TnYumngZRgOt504EFitST+wJ/krxjBpK70wC1fQRKVW
6tcUhlglKD/o1R4vE0vSkb5fBnDk1QG6rbsR6tLhz2uoSoE6NuBXKikS2IU02+oRgUgkm4ykTcZq
J4d3+2TJBiTbEB8TrylyIAwbYzjUV11RolfKMqAFjI6YFF0NqpvTOfA5gq09WmJEqcc2LyChNS5C
onYO7OC8gEFNEstkvS4Yddx4wzSqE05tEWmaCExtdsUZARQLdTLzYLSkjiJUvJXmh0GIRzgd4fe9
lh0R4uPjDz4u90bJbqRDNstOxI6iCdlXrhyuQJdcTXeVFOSn6fauLn3V41FJsuqAhe3we5vyb5mg
mIf+Iko4XqndozVa2DWKcnlOPIzy2VYvpjJl3qq0v/9DwEMQRLKMmHHz8U8XtRmr4bj8fiTOatIk
O2iZ0LhZoaBXKzkIQZfiGw3FgkVmqIvjsuNgGtLytv4eOx3IbBCOm8B+DmcVI3Qz9UTqO/j6ioQK
EGAAtdVm93JAEIfhPN81Lwn2c7drUn/SJb03rFNezWNo6H9vzwX8naNyGn4httGs8OCHSnKkQ65n
nygXkhZ3O1g5KoDXDKLAtcvxiu1AzLk2WWQG6iliPZlY1ZqzFU1mee4CcDNrg4D2QJ4NQjU5gwQU
XPbFV9j3YLxFhg1UygREuIevc90sYb95Ickoyvew+/pj/p3crJNknuNnShHOOdO4naLdDxkgTm4T
XeUpU+nFyiX4c/KdRKUy2B2tbFg0Lc9DgopwiuSGlT36+Ck3/nR5jUX9UPBKKl94/DV+EJIZbEDk
SdaII7WF6Nhc7b3Ugj5hpzxkzx5/d1xv5+7e+b8Ejo5NB1I/VftcL0HdYJONZo1bH6K7JJTLCVRR
J+ztfg80xOrfkqzs8e8LT5iPp95c9X0I7STK22vMnXuWIV8G5Xik1N9QCIHkTY97hXg/bxasmjdj
RsT6w1L0DdZBrLYCsULA4WOrjjah1OOqbe0q8E3nHPOJg0e3PfnytyADIK+jS+4d33TrJYm631Eh
q9DjCIpQjuDd7AKtaiWKP403tfoW6DyKyAyj2IpqBZ+7+ZyijqVKC7Gh/iwodBpDum7vZnQUIrGg
prmmC3WpktyL+Oj9ajpWSm1kITITcldnYwzIpy7k+s0Y4uZK/DvA6FyOFAGJ+SNb41WGNlPYiZ2G
0ZQybC0QB89kAIcoGlhtgSl2OL1Zyhk0/WV6IkrC6Qj7jKBs9GRyR9N3yRVUf4BEKn5Amzb1hYCT
3zU/yU43ZdOUwdxlvb5nJ08Ik0ePUyJJYLtzSyhonWWPw+Hr+3y5wPhTwdBZMFa97jlxU2zf5Tzh
lpVEHo/7OQTOLfUOIEtddPNNLjnKtijnBWgvIAEFJ1yvV6C8sJ/Ttqpomdx6t6aBg+74ftOGH7LK
qRqd+T7NsdZBZahrsv0afyrAHairPPPygEzRMOz6JWgzojqoCfVRm+7mlmZFP1NSZpjhIEN31Cvy
iJ+OmwRUo+k0BjvM2m0XdJDJBTdavud6KPFumpq9LZzZ3wKSjTVBt6JayNUF8ZLrouLLNOA3BaYW
7ZgxNFPJ3Tg90Lt6F39R2Pq6YzYRKm4hDKpNueIpOt8cEEjk0vTJUiBEnRhwWY0RFGNXJMRD9j9q
sihYH6rHvlb5wtLSdeHmgJzatIIOd4D6eG5rqXUsJOYZJ0GsXcn0nHFDPDYkVarHfcSxyuitRhBX
0JHtD1V64rmGgwTEX4JgbYeJJQmKda9FA/01uqJwSy56U+vab2VAh13OBl9AM15MLcIqGwcdoiod
TSQMBzDYrJWqH2Hpr3mz0varo967WVY59ziyacLMz43vp3O6JfD52Y4DlhqWA3/lBbGTjNpHdyJR
Rezq9JeANbv7oX8LGbEZrgly9o1ThLIAJp6j+8s9Zum422/9YJOh9bG0eQTnc7rgzrgmbqnOvjmL
lK7nzYQbCFBjNw8/focN4S5/5bg6t/Fd+YP0fbVlv6ApNbWk2Gavlg328KuMZlatXTVCUR6TSM1P
G2+IEDwWeOFmI7pkhBLsGy73GbNgaoYRumxtBbB0BuhhTgy7SxgwKdIev3EEP/fwUOPs5kov8NYa
fFV+zxz7Yvgwnbub5ti6a/GhxzABSIHC8qgOC4U9GVcxKa8B061TQm07DV8EBstO69nMgbALc84d
OG3/FeLiqy7HF0nwvb86VtPnNJG79CPuCzCv8ITqavn1kvtS7CziJTj2FDtYmyq9prb4q+ssfer+
Ei6O/FwC+GvhV8jO7wUJTt6YM5eqUauPrd64YPlaTGUcaDuhfHt4jwq81axfLo2BwtfJtnUMFWIU
vYbVavYR0BEp5zVOoy9b45bAnuKOHEiGF56020fOSpgugVRZNWzYYnK+KadGjfjkhAE+3KTmWNr7
dfzEviTZzwBvuItPETieygnsT6i3Rlxcp5IBDlxn+SRgYKVVnEuru5t2PmJkNfdomzostbllvjA4
4Y/dxrcw38sGsZk7wrEfCrDxP7Y/rlRBZaad5Nf98jng2vm5MbKnFidS/LJ1FN49z7gM8WufcLYE
nPNb1nAINoKFYbJTL3IfK21H9Ruwdx7H8uag8gzuHZAvixfdwkuI6xa8WNjHJjnYqJ6xK/1ZtvNZ
y8lV3SuE7GzG2UCeFbHq2T3obYElPnWgTJGeOPq0iroDEkKcCxfiFCnIlMsUu7k8FgWRok2+wfP9
UyvVvhN6jpIT5dm+uTaAqGJ2tEyge9WGtsTQcPZK3Ebft3p8bX5HEKuGB0BDuVoVndLQvuUkjp19
C8wzsi1zPm/oIzjd0E++eEIYUidzMLe70qzYQsO7Ub7wAwyG26K1xvs+ao/+nKtOgANy9ZVu4rug
fwOdwnD9ftXdrP8+waW5DDeXqIKW9TBPyKngbIhFvyY+0Uz5+fvtL3GZE3CdiVR0w5hTuUW9WWjA
zLZ+N49wJaeDOdKlWSJSX2deCPyCTM0Wu2uDn6kSYb2t6ecuUjNczRsWrZOX8NCNh8eVLpcSMg8A
Hh5NKlbu31ULnHZH8spiolMmzmU0AFN3f4ooX+x+fwqehyHpqnqRgKFr0ncRnKW2h1lwcHDHPRdS
aCxjtAQF0Cpr/Hsc+lD5JCwtUqFZIPECGkC5DhAyrnFiW9OQPVqPBml+XZoIfW6s7W+R5sOg/JLd
UvKJh2sucB/Tw7Trtwq9sL0xzOjK7pCImKZu4URiPrL0iJBf0K956fYyoOGe6rwGApyQEexGF0o2
RzoDvxCdjKBagN08kZC96xqmGyXyA6VVrAxw26Ys96CQofsTWconb90qiHQ4LDhmptJxtsDLV2zO
5AZhkn62bHy0DhHEUPxO5stP0sETnqmHk+CCf1uFO41sEEOQY3/nC+OxoI8CJPmDZPpRVEn+TSha
ndEm79tQ6x0/8LzzIKmwOXZIhJTUCA8VcJhVxdDW6ATQYgxvTv4xkAPJ4q4AFvTrqSiJJ5+MhDfb
0X7UYxaDXfg72DuxXWc8/hJlNpO6VvK7zjt655YaBYgxGh5F/0xDGf90wycP1v8ITpw9AcmBNZLL
Sldkhm3pY6eGrPBNiLWrPhvTOGTQgRSUmH+9b64HNeIrE9qJSGKkv7WLznVIx2tbzHebJUF0Cx5k
eY45kFgoLwnyDvqhTD0z26gFIG9wlvRw8RNgFV65JXwo+qBeW3C1TD/6IqrTuZPyjHkgfaO01u0/
7+Z63cV/RDhLSPvQipja1abWWqs7IrhD+8IlVxznQvO4/0jTjats1Lv7sDvZX+tHM2ZJ29lwmmiF
a2kB6l8RdINuHDfFGJs/qc5AGYHzsEOCUKI62OZplaHITelMjVq8jkE7DOtqBjC0lwCrCa9UM7sr
Vf/xwKz/tbXyvqxMROGFn/nsMQCuS3hnjXZUXAQRZUG+dFlChazEiN4qW6fWaK72OIsHiLNrcuG4
Xb/0PNUx0PO27kVO1i4uwdkexiFKoZCw7x9d/z66Nr811koFQwlRpUwS6A22tVjOc0z4naiz7i2a
BQtZAw5IJ6Lp2awhzuViz4qp/iTHwQ4cr0bK606O/8owWl6buhKGbb0oH+0z1Rm4E8U3ccPfa64D
19ufIyVGjDroszHQ9QYfpkXEYQOFzPmO4B+3QWyoeBjXn8o7knCx21FZaqlZsNOmJdVPV1yo1MTg
AHqEtT96r8Vrtr9hesrewkZWrCcPjAbP+swyWEyKyJGmXUmhVqMloOjpPaSDyOTphD7tJvOv5/Lo
DqWhXgwKTB3Dh2HuDeftQrmeM3Acj8gDQAQXZhBZ/D39X7NnuDxKfZM4HpjTej/sZ6uWIeJyom8D
8ltGApTMTIaUsQz03KeHYK0mUT+P+8PZXHjean0RJIpQhg/jA1AuVo2viapZySyRgLj+joqQy8PR
GAhTvnMImcPnn9va38ostdCvWxvxB8hJH0KiaKR/WUmlTSh7fqOP/8wrAICHDk8rJ76ttMPUvwuV
/ze/2+lPN+fKis/deAvaCD16a5LIGnybViDLo88BJWJJr/IusYl3lI4jCeF7ETL98Vse/yRz0fWa
0mvGH+ogxEAyEZlcNU+ZSuHFdt78Y7usT+U2yI368uiIEty9V6eGmxoSkhj749XZAuok2fbdDrEB
yCqfAhuMyOZRESM4OhYOwBMU09X5/0WoypIEEU8YjIynAXsftmePjn4ojXuYJaRw2IlJ1a52N5Oi
zMYlfsrOYsYfCgFbxqXqfoPMKfcT8vbxPFe/uTQ0wZkT3kvwGun0KnpRkakuU4tmdkLMYTUHTjbh
jLk+5098VDYlI9aiSOYUl6m/6gYwjKalAaiXyQQxiJqWUthXXx0bATm9SJfeGHqxshDyQjo2FboW
1+XvB75R/3zka8gaz6yT8pCkL/hLNwj20RmPhI+DaBNadsoDbxzMlKZnPqn3zibFkWGgybxUbk/V
rFvSDPLfj2Rqmk4t8Fxh1XB73uVBKLdg6Oj21G33iFS97TFxzCdmv4uMCVavvxygDNjdFZH8FCxo
a1fTwxIqBhC+oXKa2Z3+GhKqUxdEzQxj4jFl1sbMuAHsBIfKj5YXR0Eyp01RVlVXp2X7DyNdxzdL
F3gjrt5DRbuLeU1e8q6+bD22zEvjGc9wK1/GzygxQvsSwRb6moF3hnCeUPsMPDIKeFJhEpOq8BQW
fE6T9oZGnEa5iI8Sx8wkrIyjBZUHLUutANo/BBjBSUsAdfhfjxuQ0B+pRZJEG7XkQAO8yyZ+Wv80
RCpkd19UZU/AYIjAPHlbKcDsmeU8FElAy2NcZPASftPXvOJyKb7x9KsA2QVQCitnrJd/dW7IJfkN
OoY05rqOZiKJohUQCfU967hx6Pym5Tc2JwhpX7bx7hyv6YcPRdd0/xZ2y0ettkWneJTigpt4MxR9
Q16+sqxviAr33ozWoIG9QiOH057x7QoA1cY2PbqWa+QFnX27ECSIpl/ORuBJTB5WgdGMd1+0d964
h0feW92YCN+mP9vvrSAqMhHfyUqIFQrvxVbYIXqoAbttNq4Fg+scVk0+h/3vBoBARZsijr+r4OtA
CmB4yZFn0hXEbpHNZQKmf0olRjmEk7kle4d7zcHtqAtSVgWHJql5FBOFZzBl+6JuwnYRzsYRkook
2hPcVSYLej/fKkjNsxUPcs+lHHZ/+75b/+F0yQO3BOcmXmFtVnGvPKwgvciYpMqKtWPaG746RVZu
McKfOIGbt3Wv/0XtaFEvMUhiejylyplTX1XEOQ4rMUpTDJhWL0BONmQLTgpKINg6QIXqhOfuouIP
ncv3C3pvwmkUir7ivd0Iir7As5lzO+XAoB9IZQX8no9V2z1uIU5c5brWGeCXMR5FobO0sjL3TChg
U1/6SuQcGm48AHoSCS5N398O0CjM406IxEQGxVjO/5vTTLxEuDrzWCjJTkGY0D38gB9o0TPuQ6X3
TTVpBEJxS43h1ofk1mm+E0XH4pS2JlJoUBHT8s7ipDoMsrqptYEdY6uFUTuBOip+IWwY2DcxUJFC
0ZFGFre4R+NgFgtgrjiFPmPeIaKWg6pboNrgLpSfrGofHGznHRu0asQEuM2wuJD7YMFpGpxRtV/Q
3prEUI60BrjTNI8NjS6lBJzNaqBoMFSy6jR/lY0ML+Rj9aEagnsiPLvuDFBaSbg+st8rWWU20WY3
7MCy3CkGlWWDfARbOez3lYQIST5aS/qPm3Pa60Z9EE9tNSdbqhlgeIXkG++bKWI5p+K8pXW3Jbyc
gsDPUav0Z83pkY0TO3p46AZ3yCWxVg8HDR0XSa2XWWtl+RNMiWFWl72SZexRdT3n2DpkCsXCMs/B
uxtjxb7l3YJares9EPihN/ngl7yLGZE/y42epFpf45eYmvc2yzfcdqcqWolqfJB8d9qy3IOH8ajD
SwZz/k7cEyWdyzjhcUhct7WI+tXrfSLxDMcvnMapWy1EHNT8Wx228W8Pzx+pj7FyjoRP4DqoY3c7
Ld3r2nnYvdVSBNF0lQ8vQiRJwAHRlXh/5DwX/bxaUA+AkNMdO2cmSK8PusUh+lUgHm37Wy+PBUVf
S+SFlMK7oVwqhWK+DgjwwnZoY/qVHQrcsYeoKe+3XFzERHveVSqQUHKlaMRQVEx6p4DfgZ8RGvoA
ao8x5oeD4x/ZIl9JGk0PdlV/zoxUs2983x9yoxjXt8OxP7m+pZNBbBu5hINs2c80XbOy8DtOM1Jd
HcApGI//nw9Ll90eebYWv28DL0Uq6Ykvw+QWRP1FqENMbodkmjA6npgRY5x8JyH+hAi9+fQdwVYV
8wFH85P7ylaNSq/VZPqSvCIqUVEhmSvC9wydVzWNrd3Jz2S3fZviGhE5axXjcDw/3wKXvMZZdfEC
WoC/uUZYnp4D/7ezpmYDqx5NWhPhP5R61FRMte1MhPxSVI+NU2zJRrwXTnVj1yuEOijNjzeoJt6Q
zxTL39W7XA7wsqhKll403yfrg6QVppfwa9MAa4I2fKuSToxl2mwzFNaHwL2bI6S/
`pragma protect end_protected
