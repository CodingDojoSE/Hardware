// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 10:40:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A84aRQtaaE/JrnGPsMR6tSyJ9x/hSFv7TfZphkEnzXIMvq1R00eVSK7fDWzjNXQ1
SA6nzokzC7M9xdOwjN2jTgOPZyq5SpquoUuC/QhBym5Asww+JNOPy46rC2a3A3/L
HpL2QtHtUt+EtTJxJkxHDlT6h3Uc1Cx85LZT6VLyHBs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13184)
nYrDZ7nGDflsabpVPPIjgusU/AKl7R5C5DyCRG43HySSbD2jWXjoV1mdUT4QIOxW
jvMZ2+AX6eBM3iDFzpmpfwHH3y0IFjfvNexLDSwCv7Q9VCiR1wYIRxRLy7aSdpny
Ewe5tNDMB+87+NEmPGJaOnzCi0NFVqZC+DLRDN6l1+URfD/k8ZaJBZUDoWbk+pBs
t11UgGEYLvqbFcP34KtjBmG5d8cJXIr+kDEMJkXUHOEmgSYiFmOriXn+NkjKs/ln
B3nOhgK6+igPhqsTRQ1p8+HEt/ryRmZkUOVoBUTDSHKByhTdlEcKmzQbm+TBu5tq
MnBQT8WA+R3oQqfwQ2os9G33sDxHzTWw1CX34f7J3zxAMWgox5OT3B3T5Yp6fvGA
53yMXM14GubVldM2wKn4vkJRrvznYS4ftSOoehLf1/qXFY9N/OuOfFpG++2o9EHT
yN5LUGL5IAr8MSec/vccxtxvI67zZWHEtLI8eJg68ZoxR3zo0WkYGUIvy9T5nVyt
W0Lhys1BHX9/HWargzHNa5vrYlV8NK1OL8zNW+n6/O0IqF7vla/CJrEP5av6uv6z
pSatvscJj4xFgv45uJYsyfZAJpfpm05IIN2yieTRmn0eEqXmS0iLPKkSHi2sIY/K
k5c+av1PG0Ikdi8x6YxPez+vvKQPiIjO8PU2OVYnxEIU/N9ifJPTcOOmPLGJ7MKD
rCZcTzxiD1QNyeibNHIfwQ6TaoQONDi/pRTN+7NUgCVZJ/G042Ub3Dwo8K79o3Zw
ot3QedzlwAkqwVPWYEZqpKeGoUzNCYDOJG3CscTPi+qiB6C5+RiXIkV2nVxr1PuO
sNHUy7RDWlR7C+cOlStvpb8L1CRR62td5bB4BPsEmKoc/2vqLDzXaxa7Nos9OsO+
1SbOgFONq4+tJ0vad+IWbCaPUib8z1ARPcby38sWCq54fFJtKQ4EV2yx3l6gVgAf
396javurN+1Namq/KylA7ePPbu/6XyZPOieYLdkrI512ZKjHlc9ss7ncCicmrcPw
J++KC0+4CuKywA76Uf2Aw6OfCPx+flu6zwQpds39104UANUMg7HDwF/nWP1ba/KR
vHqKV+Uk+aATLNqWESJxrYJFqqhZWCdULaldQHWAUNXxQzy1L5FcJEmQrOPXVune
b9euziRvCG7MOF/uYzl68knDGRPSQVF1drjsjMpqzdA0SYlK6iqTpsMqvkV3yq2n
oMc90DVMj8VXffsQ32UPoVJcUheU48DdJ8qpnGsENG5gi2iK4LjGM7CKDjdLIQqA
sgvXELjIo/V09Q5I0kNlfaXAwy85QtDC5qZs6vW2fegLJ+6M29xspR8wsHhc78Gn
lcyXPPeFLtA+1bnyKacq931sYQ0/teuBAe0XW9wv5k5PtmdX1xNhfobPlGvSD+vy
PHG2QSFZa+SgfVvV1m3o0VQWP9zxq+JLV/cI2jpPZoA0umqeBDBBGL+lFQyp63Mk
0/WBfkw7aOIhfYcq0yyYIZX3Q23ENf9tDiuYOuqkYkAGXYVmJOMPYK+I0ugJt+np
823tkbZJb0UnB80sFXnaIxkeOhK+b1Dt2BafpjBrr1/c+BvdCsbHClTwXa+gpglf
jLGDLaNs6ZCiOohvVRzSsMiv9zA0q7suzRdNRWdB1YXLbooczzLSABsdWSU4ni3l
Tku7pFSTOQkCAUj0W+Zs5HvXlc0xTA8RdTgHGYbsAvTG5JM8bRtu9NjqObVv+8sn
V9TJegCuMARD7dUox3MN+sMUwEEyPe0p7MDTxCla4hZObLUvcd0wxByIeyqrnUrx
7uNUIFTCeuy+hq7Ulcw0msFU3/Idma8swvlyhHDC0/goIbTSaNs3tS2arpAsGuQF
CAdzrBgfX0zO8TmoBKfY2WFRV35wx8k+1D9S2lc0IYHI1Zh9Vjw3iCcPySEX1f0F
U6m5/ghZ79fg9RW6m2d8xe88lHTGRLJMmI6lf2WKahrzyZlxt7cgBkM0qEU4WwT3
n9FWPOahGs0fR8omcDZwgWfF3u/J6YPQ4NCUmr3ujNlYIEcY3pn7GnIQeaqkaFXH
v6LwTclVpbwpGrHsy1A3fEJV01zKEd3yTNnLS7gtpxXuqMaGQuiji9yuO+TTF00w
5pxySC/EUQNjT/Rq1EaWqQi8urNlWpmz8KkuXo3dInqUPdqh6q83ZTtKvgYVcqLt
QigqgIKCU21xJEn7FNskGETTEaqcJb+Ir8TX4Mgq44mwqI4gZAFhTpIFGKjbQktj
BIADVgfxk6dKsSWIZgLWLgMlN9wUJvwyc4072ozr29OKLCiCoeqlKdscRS9oShVr
aZ1Xf1/N62GChobhVjckgn+DUoEFqhdU6+OJacZXDA6TMRLir/65Ij7H4OMwyJVN
9xlK3S89DftMBWg6c2aPo8goSb4Gnpwrr3sDWXkMYFJg8/5zinb6lqikzReckCgi
HUuq2K2P77yphsFqVKXpX6gD7NKBv7N7LoYVNiyVvgsclAwN/NGFeq5rkNHR+q29
oJAEQaZw0oaqV4NRMhIBrE7qbiRs6zRaK2Ut+BrCBlVwESWlhB7atuk+5xSePCHp
lq4aao/OhHDMati9L4Dcw30sMxJtKdRdPNI4IUqU62bJarTzmRvznlCzKGybQi5k
nQyiJqmC+5pC3pV2lUz0JnsB8c20MUYD7yZWa7iOioxSlJmULmxsdO1vgwFDqEYW
b8Uu2GqwDyFLmplT63OiZZkxiIl8FsJlJjjszvfKtB54Q2+KXJF06K6x4uykGKMi
OaK/mSyE2ciDdlOE0LsZVbPduF7EFu+qqOoyEyZgZ32gOG2qpr/eG9bv0Pr4qEEt
GqI0unSsqIBatiBzZzRiZiHGMu73LKyT5owwqHxKbDvpYSjAMbPwrvYQky9zEWyf
WLncfWKrTP8pangPG3tWhJnixFbDqK3n0ipPnGwXayuEtgNHDp5+tx/eTGhAdgY7
5qWBIVHKVIrdc60oemNFY7Np6EMfOzSYLgjgs8V6H0W1lA/MFYU7YMAmHnhNSthw
2Si17QpCUzBXb9FfgPJulh8/8OovPFqZemDx4r9AQCHetlXrfLuQdyn7e0/h+V5N
gTE4iMoGGP3wZmrmRLMYrG87h70LwZYarkGL+ag/VQkqz0xswzQZm3a4ppaU3fUO
wDhVxCexAZwtmEu9W1KSistDzWkKPz1nRkK+gDQVdgJBeP+otDgYS51VsBheOJDv
CgC9RIhQQqMIpxzg5QlltiFEJw1FHwzbIi8ySKPamm+3ET5IrdNP4A+kqAOxE4BG
v65gCh36JagukDD7xCb78Yk+vlGzkv5nlsOg1VbmlBtbVTmc7VP6RaZH9QDQYqlJ
wuslCNqOJnQw716JgnVBm8+ZA8s/RbnU2AsR37nkJIwgnR3gZfsAcvYNRkPdT/zV
tIUKdqoHVgqnOGcK4c/h8rQWwG/nJFXbe6z4iiPFFtF+o0bITmsJSyrNSjTT1nJW
iQrLdNUKUAPe7NXYhKHwGLETTepdvCliJnhlEWIcFXRbgO6zXLCJtZQ3DbLSPh+s
t4PP3IW/vzx6lTHX+cyofDEiH43l/lTosSuwufJMlRodaJi33201JH41TE9E6jWo
ObdBBrdCzhctWZBujtpphou8LLLd4K1TTJR4aidHerbJcXEHUKGVvc56oTQVmOUp
iC096WhmcIsOlPKLr/Q9htIIS64YtFdIY/2NoZEc4FCGM2ghVelsz/CFZ7Ij8qL/
3DvYH2nhW/m+BlodrxqyHnKYXrGiUQuHXvXC0hzI7mBsix7JwbuMc7iWgOCrgjE7
0oTf/htLmb4ms0VrBJe6Rs14eNqP8RP4DU1PVq6AwyZ5k/Mx77Oggx6CrtxE97dQ
FhH6kgJKX2TZ94iENqlTUAcrx3MTZQkmx1kxT2QT2H0rid5+Dnyk21eTAfx3LDkK
cOu50g/0BEyg8Gh0upGb1pt0AQv38vzM77CELyOh1Rq73M7dN0SKDQqDVhAabbf5
ibV56HxqXm+HCqZqMznZNvApSZURg+6+bKGdOEvOD5zTufhWnH5nOW6vER2caJku
BO/Vi74Az/fWgleDft/n0pcRVN+tIrJOCRhjW6Dsh8vIzIG3JJLq++jd4tMwFQ6m
6ruipR66AHyX9BC69xNwAwMorR3IJfEMaxDoUG1seb3F27ifq2S3gT1YkH18JH/6
5tKlYILvrLMrarUaB5yP0Xdbg7JNNG1dxMLJummPZB0tYsWQ4z1m9sYtU7UtPDCy
7A8dW/Quz6yBy7knQcANi3NKq2liStb9GMzIHi20zQSgZ0j5OOnkrYpd4eFqFLnE
b4Ctb2C2hfUFmh48UXg9jPeZcomUfW15W2BA0X1L8dvahwlcmjojjZlRlcuy08VZ
Jzmoq46fsn7S9sm6+aj7b4nx+YR1hNhdQjN7+8AL2JJ/9ic533QyhasneuoPYZny
7qbpvEvOXYHW2wvZWGuZAQc18bIJQYd+xDKJ0egko+qcuMuyAQhOBMOf8XQg9R6U
BUHD7sek0K4lwpXb63JxTZsUg18gz8i20gGbf5BWr4vUdTWxZLuZZ7tpRYugXCfY
qzK/Zjlq62gCNclR+IfCLNdwp18PPPXyjYcwZUiG2+D9/BfzkxLir2sWcj28njQB
vFRQR72GIW3Lgdkxi3xTy9jfjdJI5k7Wo3iY+NNfKBoeZH9FXjr2CPnaFnwQRNk/
Xnv46AWbdQztTq2AHV7xy6YcQ1/WpZhxISjkOnvIA4q9FO/bHYBubWHPoZseFAm8
90a3ZJomKI+vB5c3xxDQ4UQkaPZXaBjxYeNCh0hI4QJMrwPGPa8UwH2vV8pQu6/P
s7Qq0sX2KgowGFYmHtMSfCL+I5iqo1VxrqplTYeZuHpoPFEu1PNGLjRdcyFCo7c3
L0f9ngKXhyLGyV3FZpmWkO+yjW5wwtjWrmlhHyy6KqTeZe1uM9taYWsnRdfFrPQc
EkM5ijyE7XatBOJKE+PV4w5seKt98U4waG2gyBWt/5gmvqsXjB5SMZqMgiM/0kCM
BaXTZbSZckstJt/30u8Fenf0hV9w0ApEsSlGJpg47UTZgThWZID+GK6IzOHQcAw8
6dga9DWY+m55ZHm1E8IUtbFIOdQX2c8kQDNNWkqwO5Joox6mTkhetUpiOldi0N0l
7cr+7jrkdujINO0qEU8wm6M6s7W50c0aIQSu4atghLZTErgPKDfrNdEY0e8bTbbL
ewb8KF0aox5bZpyu2IeUrJOFI9zZt5KG+9oaVACpUC6K9qz2/pOYKmoMbn7qCGb+
xn2rbq8XXlKn95NwoBrKd5MJ82QuaNHN2pVb+7PbQWt3vfSjokHStpgaFPYgbiAm
1D7HpOMy1LGZcJ7QwWyg7tVcVvgHZg2ZcCB8p1sPEYOt30H2sRbix5+z1Bm5mpy/
uDqWaNCnj5FQWwcD2E8cuD9V7yjcaeH7eq5bwXh0N0wfECy4K5VuTsb2rArdesDk
gDqUrrDaG5dbMXOPP9DOGWXIHJN/zvwXja0rkoEGE3me+jONxtX6Gong9fyOMT8V
/wb2x7PkxGDTjDF3kL87Ecj0b820vfxWT2jvYvBxPCWch2BBTiCTHPlgL2i4Eskt
yGaXVwjlHQVNhxadUOA3RRUBCnlcyh8TM9h2ynfEBrsCIX6Wmowi1ootp4/EUluc
pijqG4W3jTGlvKXhvnDCGiyv/TjyiUXTXEKbP3kV8yC3bOGcEDFmlwFjqmazhXVO
VWg4wHY2NPXlkhCZPOLjOQNJ71Fi71NG4sPT+JfyiPLM5y+Og1g2m/8kxiY2VHLZ
Ik9cnKraQZ5w9ka30XVclQWwE/6uj6+SutJUWv/LdHP123XElOkDezyIgFNwC+9M
Efz8r5PGIC/nK2SRjxjJUqUVPxEO1nwg9CpdexJOCdf+tE6GQbihrSR0fiiotBa8
vCDWjwYRDHPY3Ae38Ly/G5/TiT4DXomT47cT5bPViEH33e8WzVbURt1jBj0LUVsY
ao5j7p/rVRVFaySAnTPqCAvnQAyyWDwrPxhvtKHcgYgSXLXyfmpIS0rT97rfVEKw
6Ffaqe6al6+PNkpjR082OzZWQqBYhFlgDb/Zm+KpGH57OdvgRa+OkJf7QnRpxm5n
5QVgnQnqbCiySylbGV0hMKhSbpirFQMkdJXVqgboV7/QsoD8uHmKlPzRmuug6Lbf
GNL5WjLlg4bMWGkoXRxlLL4oZCm0NA4LeXrDSohpMom0+9K8aTWfBqdrW1IWvf2P
4gfbcP/zHRKWDPvsD9nf4VFVtSCKF67OcmKN4icbSG4M56oB/7SpAgnhqQ8/nxHS
8yOgZpDmulZGnKX4P7lJshNHFnTaa79hBKcXSQvIxtu2KbnQQAjj6I/CfAm2z5El
2roPvvJmN/fkFeKtJbyQ0IibTZsuDU955vq4M01htY2LjnaxPOTlnq5tkun8xB1h
xCxDHHIEE51GxwZahlUZkIS7+WNp5rqIUYjYaGYXQFJfWe2i2HWehcvS/37vkaae
OsSRMp8KLLi4xZa58IIetvm9yOR6/ROWMgpyrC8OsxJREBQD/nzfayRitkmJITLb
OrJIw+dUEZ6p1og0doo4hoK0qeBzvy/pJIIZ0T1GuQCSvBdEaIFKE/eAOPdHtNhz
IwiIvhvORILmKsUBhBfn/tKslIgpOUb46KUFcugTstQf9VIzrEnOmtgufk3tWYp2
rUvw9VkREfs+1ogXx6tdioBta2BTUdcdhRsGqmWD99XTux0pGX+4+nHf5s5IVINK
bH7heelqBB8qkzN9wpU3F68YiXvJm1r3EXlaSqRcyq7HNaMIW9J/Lfhyq+hyKzYi
ZF1BCXtBqisFrJeTmnUQuhg9ExA6yyg+aC2q7m2zKqOqga74FxWE2XPlT0gSigyM
PehEL3JcxBGqvWdsSMAXJkQCRGWNF9n7FP2lj56RUSbObi/ZIvi+7W2HPWbzEqZ5
TDZwCE/efeKRjvn8wO4vYCGbF14en11SRI5RIZExgwYndgoCqnGTxU05aNYNPAkF
0xXZ3fX+St2vwhGhswRgYXOFAonISabTspLTxpToX4mjCIaUsvyq2gCTRrqZ2pRf
iJfpVoRW0S4MI55j1psOKrtTQQsD1f3Qn0G/QuHSP0DYD3qNFbKE9LR635kHkUF+
LURqSRM/BH0vE1cOZbNY43xR0MC1Z1pGA748uLVnI5e5+Ax36o4EpAfGbMvPEEIf
ClvAQQxNagIZZtj95TGXANe3pKZcQdv1N7dr+ttWdVMjTIonceC329RguKrxXqTz
/fCFWJ3z2yFkl+9H5l6UEwqFHgoWM2QPsQstWJJo9aVtFhl29BRbwScf11p66hnO
ZzterwiLxKndIu3mcoaEI7HhHEr0pdAQqwMvAnH6n5OdFit5hpbxJclGzlgCR5KM
948TTzCr01dGhb53BB6Sry8MURmWFPbDY7f6fqj1VlbKyMXYWvjoZ5wliNP+EYt2
AtZ4tlFpxssNxqDVPlBRKeUkmGYSpvyoq+NUTeJAT41jkylXMxtzGe8Mh1jSIcGI
EKMRZvoro/J5egAFc1QQHza2K/iVJLcWlXJM7zTUUrP63IhlBKcJpINcJGDPCFpA
yxQlrJW4oKxGNWMZtqjcBxzU27KI15tKaZvUWqwMo8L+lojy8xGXPiBYxUjfyk6y
3eXlQWObzbKz/4KKqv80nWkfEM2ktB1q9iSSDszuI5vrA27pddjPx3oP3Mlcfy0z
Mmj2kgg6jBa/Q97w+JlEkE17/i7P2zjLY9d/MrsfP0VN+AJOENJK4Xz7i67NkFy9
1u5/afzoghVRwefGy3ltLcjTcgi7tJDVcnr2WJLrfxPxd1OClWg54ghHjVIKmfjH
xiH4G/e2r+xHnmS3Z71I7A3p8OhU/GJwwBbROrzfarxqCUQJl9a7isXAmw1RjNuZ
SxF5surA1Rex3X5hbC5mOZObv44XhF9OIz6qoumTmnSC5zLDBLm/zK8hMSCw9zNj
xyrFA2algZG43dTRlDU6D90cyV5NXEIoRe3UbsHO4VMwMAzPMJLp2D4HPzh7wMhS
c4PNTyitmi3R8aMtt6p5yMwxnziVZZECbJwrYUdPuJ2kvAyOXONeIGmWe/bWO6ND
YZBB9UF17tm6YO17uYhnk3toLD7UbWIFYw7f7AEGPBDSIBFPAD2XK5vQtlshF8PK
qaImxhgEEe2ZI+prvlvkgPSs7vdgCpttxTuj+qSscF1XiQ0SKXGgh5A1+9p8IjNR
jdcpvJ1sDY9EZy69pW8YRzx9DMPVpwMwNA0SCCLLihYsfCur3VXdA+oSJw1m72mQ
Q4tHXqrkMetGBcAcS2/zzBdC7ZQa9SGe9SzjdrTZL/zUvxA2AQf8j+VWYMUgqpSm
MG7RhFwJiVdFpm572ckGTx7nDRF1L1/A37gyZdxvS0NWV8ZFay0DkxssfhMfADw8
7pqHwZ+1ksZIgwafSpwk1THe5VC4HJAlgP3IMCv6IzP6Ld1eWMiKBqwlqzJLZIu1
cUru/qedYW/Rl8yw4M7Y3NlpVvRsj+/RDtZccEWiKdYs2bXxDFMYPCBOyWW16vAg
AfGbBEHKqqNeqiSLnj4JBItodJOnpFJhSc9Mg437KoVHFi7VBM3/V/b1cwx+B6Vg
Pli+1Zm77OnJgBobFlJ46BbprxFWO9F4axNpT902ETJgA1nTUl/vKw2baxFBfhl6
CJ8dMBWYGzFImZ0C7Y2oldG7nWLAsZqXQep9Y4q4glCIa1aJTTfwvab+PLDX9Z/+
kE8ONtf/wCsPpOLgOECazCL3UrLICPFVCiDll0uL+XLgR+7NErUXowRAtcO86yIi
Ai0GccAz4jO6Zf9aDfQwmVVvzXhXT5WYUMAVsPKVtdEiVcq4mJb6haRSJBY+BCBE
S1ZohzzvlEELWFjwKmEhBLGBGBx5Dci0lAT30EzugRjLUspdDv++x2dhQSG7Ao0X
HDOxram9algrRg7yInruZHUqV4hLf7ELqdNhNk3dkZ9VNVHbdG2WI59RDBMnP310
iW/XttNxKfSh50n+5GwnmT5PdfRijVL0CL/9i1HUlx3eLLGmxN5CKMR7pBv6F9em
CaDRqtB8wbboYIf0dAM0nTzYN41acYX4eQmlbp40P+w80ndt7RdD5CWHSfHXasH7
6Wi9jBAUo07qpVaXOWKcBtr4m7znml5WgQY5+gNguooeuJxrqhREGMJhdjLkr4Qj
gnUD0JiMZiefcKyncZDnCYk4sl/THuxxd7YzT2G9/Uq3RjjWmxoukx5J84Cwhvom
20eK1nnBJCYO1SxBtYhptv1dGSwmCo8fNhALtvJxzXIgplvjS8+e/ryz1x2bHGq8
gtUBan0g1d0H4W4VqLkCX/qx9qfcLwIz20teQKf+dOfkbLhRipNyksidYjQUw89Q
yR15YSvYMjcXSHjhblojg2fteVIUj8pfAl8nRHsZ9h94L1RjlHgkVGVWwIzaASQ4
EpeVQKcrBlAsGpJI3GjagUFehcZkmX++9embBll1xdcBfO/UPt5K3dZUplFc+6iW
3wzVzsyE/BPSTItxKQ93GSQeBJVh9SRUCriIckno8Xjils1OFTn+lFtU8m8ub3H4
4WQJKlDVawxjXKwhRxZJu1T+pFUGYwORgOLO/qfTp/AaDDdt43ncQwX0HnNVPdXV
nY60YdBRduO1r6BJ3UHyerOEWSzYTPKjE72PGjH/7XsAfgb8ppscii6wzAOV+rVP
bxcN6M22oP7lF5q9HIZKwbovarvl/8yc88WAPNui1OrNomyNzFJFoUcHqebj3Mc0
/4Wo8sOKgQrk8l3/w2oW0uISy0gn1apcYg7uWikOTYRO5S+X8BTPUyklfny8be1/
YVyG3iZ58Uq8ySPq93TOOS/A7MLarrYmG75e5H7kSu3dA+qb0pfuspq+RU05e7GI
z9gYm3DiiJrma1aPQX+ZNZSgpQKV0AXyVUfMTctLRwGeRZthX+9OxM76Jl61teT9
+IKhE6+vAfotuIgapIJc95MEJQzVfs6tGPbZ373tLYy1k21WqYlV1AP14pENxTY9
8WFMikqrj45tyoXQ2Zv2f8iy0sn+6Douw+Re1W5ZswbV4d8Lh0CXQ7ECMwl33Ror
RI1JTtfKKnsbxdlnTbLpV/KafG1kQwjDy8b+YxI6ZcVp15HDKcFXIOwMeIlR1Ps8
6vtROhxakPP8SvCXRFn7s40y6NR3PQHFW7bIAp1l2VcCUXikrW8uvBFazsZhIg0U
QFkjZ9I2lGcit4PO1F+vgWX7l+Arp/HIm7TF/15g9yv9odbPaLyohAKE3wdHJG9l
+PW4JkK50AvPxNPjp0fBPimBL5MlUsUYG1YbM+7BY4eLg7/r+eM5r1csac42B83p
WjfDH93K1tEUD5SOHEYAg5EWXLQqvz/qE87VIjFENUtSJC8n19updbkIKnWL8bcc
EDXk7S7uh66VJPJUScYv351x8FxWbTzla7fEgmRRaOGXXW8e3vIE9jzNaj634Yws
CO2S0thQApU6zqzRjcfWrhCI92Z9GbG7AGz6chmJwIidQpI8YoCYxnrAeOtNcpP1
rWMHrqFcnRp8LRMP9nPa5YEzMmeonf2/4EaYDyuJLw8qf2r5X662YgplIvkgruU5
cQ4rmghxgl5mccBa38NHxw2JPAPbQAJaiSQrIxHjWHsmkmRIM0FiPUfXJs0C02hy
tTUbEvWmmh90zmaW9i5KcktRr9yvkUqIB6zQH82MjoAmshyXN+wcaZZvoYL4jJSK
oZZgDaZ3cNRM+KVsd/QDksNto8UpQD5QcpYuTnDW5tPfDZXo4Dd2/Av8Pj7vHHEZ
9SjteP9AlAFeDCMEeX2RVNEaHjWTy1ZvXEsuS+I8lN0cxnpj1Ze82Fs4kSfSid87
IIa3obSE3SdK4/oP0XjR8tV9rAgOWGFKTm1h2TDHBd4RrgtzDXMhn1tpKBOnKfO1
x+dMvmDCiDZ76mikvPBBebZYetYP9eYybgRLyaJveyuOj7qyHdVOsi2q/bLwK4+Y
o7i2bFKo2efIckgqPl1KLkujfsYhZDH45R8Fjhly5hjz/RnsXB2oRi8LXv8Dheie
U+w7N+4rAZaIWxsSp57n3KC98WWJKY6IK2BZUDhGxhWwpznCXcS4Mp6t6UmtXL3M
5piQC35y+ZEgSzhn6qqfUJPPU3JQZXcPawbKObrqPNYgzVHGJfEE51mcfQhSVnA2
jOOsAMxY+lOtL60dFemYtaaRaKv5vXHS4z4WAq4jk+N3CMBlpZZrLNkNfPwTaF1Z
JCnvxT8Po2dFvZk9kv3I3EFD6g5M9FQ/bqgBgsGze5GySVgoGs84Ny6cam389SbX
uHkroqP3sTibusH1RGg16MSP7EwIalokhiV4sLHiZCS8eZYvb20PJjukOi4ZMFTP
2lW+NVR7YDmCmd/BzgAxCOG5keb+Yi/GpM0IXrOyghoTg1+0r0SQdd6uaTYuRXXF
RmwpIaxwd5vg3U5zvRa3LJhoDlY56I44wFzcRypd09JMUjThCMV5RpzEtmzduArN
qrDAVMesTHoGWb0iwxuKLstsMW6H+5Mf8exkJd/LFMRqlEMsQrUxA2ox0j5FBDeB
fZvKR0oQx78CaNt63xj9CKeB3KTO4sKoCmk8J7DdhbSZuVW0w83fq1H7WXDHNv1i
nPL4CK4JEoYQG3iHlshEeoLZnrVysRi1AtGohGmMsbVeYWrZS2xBXuVBIba65tyF
eW1dt5+WH5apz4AuTYcv05ZVBfnKQ/2NK/kmTxlHT2TZHMkBJRZfb5gnu8qoR5y6
0WLRGiwoE2TN8V9ePTV35JzVO2ufyPAXp8JTwUhgPLWmgWvp5HVAUejYVRuDIY69
qJ5qBwK/hUT8mvH2JDp3Uo4tcCJhgsyyzBT4fZ1qrTKFDcsmFcs3banRsWyvRjcM
iPkb2CCobHc8QRBmF4lCs2D8i6nfJEQRqJ25hcPGHa1dgVO0eJ0T+/6r+pGDTrvV
k1uLpxg4HXf2HMUOAX+vBQDxUURrnx1YnzOAC1pOG5AJLqpskxW3Dziv4XcVk02t
pzjtfGwqwfNse7dOmhnFOPf0eInMSBFfUZLU4vQmWoDiG5Z8/6ypnKwqO1nkMmBT
n/4hibC8de8ErUANiLG0+Oi7LkiMMULlaNZQuUbMKqLuDXoF0FuMTRdCNtHBpQYB
DKgbRJPrplhypPiKZZdJXoDKis6XeWPAJwqmh94zn5rPLhuP69PXNE+N22MJX2Qe
I633nrXrNPPDmHgHjvX7dFnMgwvbQ8O0476EQT8sd+ABJeW5ZY0hV3c6PLzcLTql
HiX/p6s7Tr9QS+FcbSoNErhttEGrl7LOLwC/p+MwRySKqWtDuLl782H+yI7q+ts7
5jKHodrG0BAJr+qMA3S5n34MKvXC3T9FyWPT/J+QPUF5sHQsXLRkT1A47AloA9w6
i6/yp1VuycDyaO7vMKQIdRCQA0p8rhZ+djqKIW/EEjRpDZvrJgM9vHR+oTGiFH4/
FwioCTyCh9Qu6ZXwQnj9UvvVDhuBzJiFJQVgiEjmF+f18CkANm3tec9bDeFT8nN3
mMU7BTUWef/ihZ23kBJVM9MyD64pzr+zmED9TxVQVkqWwM1STOhXb41yZM7GPcPj
Sa5Dd1FG/6GktmpMUW38J4rtNa4a2GIO/xxqHg86xFnuBynYtVTMkXZ5lIjEvM0k
+dCVWpzXwPSlgBOFOfezT+v+OJRQ3T0AgEM/K0TWtnhAe433avM5P5RRiSRS0zau
Yg1zTHQlbZhjARa6n9LcZVFMTAoJj/T9zT5Nf21rltAp0U8Nixve1f7NwWj3x79H
QKkU6mCWUlZ7PMMJAPv6ztkb79V6MgjTtcw102E2MnjqTmYn3K/N+jqYyriu2rVg
AEaRiLldGTrYkPhnh94UgeYWMVZWzR+tsROuEIo2h0YX5Ewo5uJuBDVWNAWgBiUc
0wvGsxj25I1/3lje03/KpML4XLZkkBiwWuKU2+w2cswSjVhqRfgGbbLrlOPRCJex
TjuPIZIpIJCYmEeuzVvBjWoYh7KDov5czWbMa51roJahZpUMCzXmnsuJNtIaOJ/7
mh4Kmc2tyHf62Cz23AuOztSq6M8IUWKmRz/Uokkh7FJYU/jSOqSiZj2BcHa1URqk
D3wjm3sM4XCoGoAQ8tbM/4lMTWXuWeH5pqvJSmST2Zu1X9Sddfup3RVdqFDrrzGc
21SaXcAPxUaG5RDF8KmQRotMtsvO5qkKnXdrXRYCBCn6pXlKyJAJffYHQimZhTo0
fLKetRfVYt5aCLHhbVP1iWW6qqqBaLR3freFXGbPc6qn0Vb9PICpvZGfMn4/BPCQ
mZA0LUXTF3udwhpAFBkkM6xCJyXv0CplK6DQc/8R0NYIWswzgyKQKZU6/KgpgrcF
m5qkc9+7odag2X2m4jQmGCWx6wsN/gWYPXo9FNZsSM6cVd0fddEPnNfapPn+xT5S
M22vywbSCUOBa0JKU433FADAOzXlgVnCELhOrBSpM2LZ92+Ty19FRR8r44bkvc/P
rp/eK1wdq2+Jk88pOYylM6ru1N4Hw+LIoJU5vvRfoAbf2B+/PmOnDJF0UD4uJTie
saaVW3+d7pCXVfHgvpu6xZiunQtYdRdUk5DZpbFSNZZtYRS44tuMYyfj16tchZF1
gOBzC1Q8Ru1FGf/eB6ws1qIzyCP9c56E0AH4NxfdUL9Fc+nrn4l7kvRkhHZYgN2f
zuyfjXvNp/63yDUNYXdksgRGHmTyv8Fq5RQu17Wd4c6ABNyfUmrEhPu1Cttx9/zT
SNyebyy8sTVvq6PTe+QwmTrZURm+NtqHSNCOWr/Vnxd0LTvRMureeVM6Nkb57Teo
lBBtmrdGYlyPPjCtCzjLQnHKMYljOLEKfm6/1FIr00tu4lFpJ/ttzWqr0HuHXF14
Ka0+8WMUcXhubXEdhFqUdxuzNEbnE1wObuYHd9HHatSTRMhWxIW7ZKwBnnRObZ5I
G7JxWz28Ga+A3mp95TrDi77c45bMb/tMsQsfIFRs9RhrOEDHs27BF2QoLf2ni3aX
tljIONg4K4kYdPqhSrTX32JEIbdhrdeKq03gtFhjkGlnq2pOV6wF52Jl1O26izsi
fWLggJDUE9SPvN5CFROD2+6H7be+8q5+s+9A1TwoSVR0gIE99JfmpDusdN8/p4p+
vdr/g5EAaCCqlg8vexWHtBeBseB1/3lgECTJMEfJ1THA49IfMkMNVeAvVnb7WBSS
rYhyeALU7It9dfO2+T8RGnBy1WWgpSqKY1Ui48CGlrG6Sh8EoaDFvtcFu4IOaSol
vD4LZmyrHgMC88C7Q546UIxGXoeVc6+Q5aQOabDW3ALQjym4czdZLtPkOHwhmKGA
EWkhu3HgxjzdLbfZffiOd70tFkbJzAUN4KVx9BMQpHljscZscgIs3e+4Swt/93cI
K8kpDXn+WSqaBmuI4iUBqNQIwy8+hozvZ0hq90p9TJTXmEvk+98CvsCttfcp90gD
TSgCifGtny7oiAvy07OoyV1LcIP+05Dpe7sV6NjXX2n9jG3rg8TtxUtPHt03HYgU
2E1O1gRzck/tshR4e1OPf2/nhc1RPpohhRr1kSJD/XKUOQugrfTLa5qPiEaRDGhZ
7sLMHfzBP76nR0KvEab8hIkZ88nZII1tgyZsP9zlE9QE8iXrIwSuDOi/EmFjwD2O
KHCWEbh47w0rjtshJWrlgvc6GFDIq4LE9cNc8h7rdFwP6f2cFPqXKdcd9umU+Rt0
VY8XY6BhsiGfQyk1Ufnq12tix3+8HHMfXtqvirIA30eS4bgLgCSGMYEbSfIlJ0mz
eO9+lNf/3OXxOBh80P7v5J8xBkfYQzenrpMjwEgs0S6iqhfZFYbs0x2XNJgOb9Fg
OLP1iyROMDh8Lz9l3Jb8NOkETdm5oH4N5ao3zwVRQIg/UNkfNv+aEvteBS5QBHQi
x/D5+seHyBLFhc3OYKamlpQ3gqf44PESCr0YOUGZ1s9lrp4SUVagXFMoKCHo2Wi4
PJMNz7MFMAn+8b7DoFkFt56SbI6mTuDrc375FDZX8uJuvjkcTlYam9sPsxfZuyAp
qBwhaAeCv1i0riFvgciiJQCMaJY01yn8tpWzbsXPy70Qxj7PlDtpf4n1uj8uPHM0
SBtq1N6sMoV0Lxq5nSTH8I4R2uH0kBz9pVt6cxZb4741V52o1jqvlo7xkxvTKA5h
5l5a2oGcCDMpWcCkK8Wt2EApiiGeZTKQ6IxyaE91KGdx+qUGjCJQMv81WPQpVguZ
iFLbNiWAHJRcCDfrKVTcFSlLfqJpuzz6DXQ8Gz3P26a7KLCsKUuJ3vQUoeN86qc8
7aopdhtzLu55xPasIUPD39Q440tOEde0BFUPuy4VtK0d1VhsoKHEL8WcARs9K4F8
STI56DeSIenW76SQwrmf+j+IocTiyqbhG8JfZKbiIde4imkO+so9WMtbwtoYUewH
XCFk+7n6i533ye5umSecTwPiPxGDGuGgNLrZas0LDq/1eNc1SGeGPZHB/iH5u1Ay
1y6SUrnzDIi4gX9MYjiObq2xu+v4fxWVcF8mh9Hc9387Dg1tthOietlmkKtrfMQo
U+RjNgWgzFz731kAXH5ikYfxuvwawJt2PRxdTKRyZ5xeEcSJbHmSX0u7A7VBdPHc
pTyZx1ds6KPIFHyEnzIWbj8gRL+cz7rsNsp8e1bJK0K82mgcpgUvVCmyujY/JxZ0
wbXSyA6coCfVmFrvwIQpgSYxZYxSwFWjLrdR7Ro2aP4LP26bLLdaQIAmj0z9VCrj
YugBY0nFaaIK9kQzZUjdfyLVz8TCi/qvLOqYzEONUeduXP6oK+GiBvU/WGwz43gm
caARozeeiZi8K0CBgeFwvzzqG9OAtr+f/b8lA+JxwMMq4li6Rqn3J43hokOnvOI7
21e7lxSPMcRNevWTriWFZJ38ODl2Fs22eJGUlUhHmLgHKHF8Sg1xdH6R6mCkktu3
a7eKVrsND5RKhNKYnODjrQ7FpwF9AfmfTCEKucla0u6nIQal5l9UOT79pE54V5js
hrw44un7VgMJDUfPD9qCxIt9BJj8oPRdztgsRqnqdJs3WsUqL6IriIPLwjIB4mWo
juWj6CUUjroUU/aQsqXdlJyHUMhn7UkOkd1P5FxEPo2tU7OmQ8kVbk8c1360FOPC
JEgL3RV9mehZezqEIDvj8yzsNuGJsCObxX0XGWRXp2AeGivc2upGYpdCiahK8RfN
HfqWzzVPHwOS9WLA2ocntLrjTBabaRV2bIRH+etOuLwQ/FHdJCgfm1t2DHoAb4JZ
AEecO/82QkCRltl5uWXD/bUaelgzbKuWMS8q0Hq86qgUtobnsfjI0t03qqeeJEPt
1C0LAXDJ6IzkrYEOZw7R6jgLhNBPpBZHKuldVfvJvitkOXXc19muyLZs2jqgmSA+
Wcld7785Gs3xvTpUSMk5S1yZbeLC6s1I/ilqiTrWcbMXf83Fkqz3XdR13+Uu1twP
KXQnOko+ra9z1BoKfAikWYS6dDdQJnqm7gw8PCmCzyMVANRxbfiKZSyrsE+HAJ0u
3GhuthbqUiu6CYrcqYUZ11V7qDoDcYTXU4MGqBqxo880dpTaFPtUhGxKAtKDgxSB
vwF91Wtf6TPe8sqnaqCS6sZEqPvpwQn4rBZOjAZT+fouuFapS/tCkpqCjZnDLrG5
DXGIfsUDqVVbxQFXOzKNZVGmklzQkw11ddL9YXrkj2lLBq9tsF/A7G60xJF/Btx3
wEbv8cI8yowJDLge5lxiEV5ARNmiH/SIsAtxG5v5dLFntdbcUV2rAkfaLnV1PvMA
Ew8gXEpcsY2nSvuP0vq8yTRaVrDYQjIu6cng5Im+fJx+0PHJLiLCCgPv9a1ifWmA
Xb1nTWcrYWAim6OY09aTKJhdiFGMUrOq+wY6w368INhWxyZRZeJiaeJbImy+fct/
P/PNHY8AwfGjNOAVy+olVRMTB3omNVUWrGWKpSC4DHQ+NiWYsD7Uy/6MzNAVqVEk
51MNOsh816ahhMupNh+YDnOmzwVqph1e0b1uQcTfuVbgINMxw7Eqzo1LoSH7Pt79
EsMkKkJ58cqX9iCApFOSSVeI5tA5+z0x561DkwEBglTBdx2qp+RxqmkCt9qHZecl
TqE62JTkWzWTbnQ7atNYmc3oywSl+yU6HYSpDe9QojpuYrkSF2eR3RIzMUJcPhst
Bqwg9O4dMcOXSbl5eMRsAhCo/RBVnuF+Ohw/7TxdrLEkFIhE1NnkI6j9IWoNF4Xm
Lpjo5SX5FsiIvuXX2gTdryrdouLrFkdGBSXYVd6/vZCpvA7ElH1AYRAUCEBVAvh5
4NU1rmdQqJbZ9Ms9XG9FuUcAMeHLJ+AeL5AbFm8CvYn1eWf8YfRXONBoo/dPGDEj
pNi3MKYIrBBTBWxO70ERqY6+PjsANhJnkuGeniWdT4764BcrhprhgQVF+dAL8R12
s0NVlK6EpM4ST2yPyT7j3KuNAAyq4GkDE+i50p8ymdPBLAu58DPMYtDWrfVwMW+T
lgbz3UJpfUlhJCsEjYLkpwQQ+OtAc06K7d/kpZ0n6BZ1aQkxWsLZB4HuQS1bNH+O
YxCP5bs9RE4dj3nswq0ChSZTJAPUBOxm5snsm2wGaLgsEw7QwWVL/Uu2si16hzXg
Uc6ODCFVSINkyxJz0vRofkxOb5oj7un4h3ProNwI+4M=
`pragma protect end_protected
