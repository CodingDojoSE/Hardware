// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H9MYYL"7;LT=HZD91(ZI?84+'6JIM#I,&#)W'3L[*V27Q&>66HO=EVP  
H_WYQ(_,8167Y&YT+C!HNH2DG=GG!^GB.G%7Y05,PW<!^-0!L:4[/)@  
HTVET.UD('J.T^> XHW*,Z' >UN[R^ G2FHV&F-ORDAW!@"<'NCB7;P  
H:0]U, 09MTA%J=UJQWM1H6V&<60S(@<>FG_L(JP3*7.^>^7PXSN^*@  
H7M](,R"IY* 4. O#H_^D!9K8S^9(\@+)W-Y4%<^"*5IL\?&B#58G(   
`pragma protect encoding=(enctype="uuencode",bytes=17520       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@ .,B\T.TM@U]E',X:O,>1NV]VTJ@9;#E2?MJ$]<6N9T 
@S5Q*OK=WR$-[(_G3U1#&/87#7TS\&E-J"ET,,CAE(.( 
@G?7PZV_2 -A8P5!!6I:7N'F%;85(X '+("W?V_8:[<P 
@=\BR5-4*P/M8RPV+GUG3Q!*5K'UWB7ZEA:D5%^.@,\( 
@-V!3#EH@+?]K<3HY?C0+3K[7,#*G61>4#YFR1E*+=3P 
@NY"/4C:P?2(+B&B"#E+R;I#"KP#H^%Z1O:*8ZLK;K!, 
@=Q'"]K_CIWWH?F0='<:Z_HHQWD=D=J9IT.^3Q*SJR"@ 
@Y4+&,+4.XK$$OWD?GB)Q'+XX2Y.,&6I^;X#+T(QK;'( 
@BZ(ISF2>PTFN"I>O7X9.*X6*+)D#6O<XM8E/=)6</(P 
@7;ZXH[VP<JCI1,HE2RXA?4DD'*N23IQPF3[A<%1[:!$ 
@1E_C^:9'$5,_\;MR^1[PT)$97RNV==3U _-C=Z_H-?X 
@"TCIX*-HR=Z?^>^^WT!=3B^!M%4W]YKW%UK3AC>'>>X 
@Z""F]$$?CS7R))LU<,/G?=TRH#AMQ-(3!"K37-GS#W, 
@^I3/O$XI&:Y8<7350P)[\&:A_CO)I)9ITFLMB<9SRB$ 
@!.M4D4%92'[!F@RR!_<^^%Z[UT>(AV'VIL']8$4%_%\ 
@"T28A <E!\OI%,@MD]WP]3/0)48925?R\Q3C1B2%I9H 
@6<J#TX:%J*G8MH0MI2MZ[^\8;P\5&1$*Y9T?E,[OB($ 
@8C+%ZXUHTE(H."$/EN_"?,P9]&Z($;I'<7(<TR?0-<  
@U8\AH:'_#N70XZBPBQ$5:I_W;?7VK0[VN%V4Q9U P:@ 
@I8I(5!X$UXG,M@>:2W>#X6)$,E"BUOD#)4[^;9S*8LT 
@[2P,[K%_SL-C;2$VG_V*ZEQ) 1M)\GLP<6I!_,0S);L 
@-@E0OM?+\*/8>\_GUT"@4[92G<JAJ?H .@XIP-*^*ZL 
@;K^6 'C2(MM^L:C+2"EO/GI#OI"&M#TH6R>E$[0LN7< 
@V2QHT-%K#?:A-A*^B./U/C>M5""/\&FTI;[ZM?&]<&X 
@E3I=WXVO]!&] Y:Z<NK>1DR<PU_(BGF$:HZ+E!LNL#H 
@%96 ,NY"^+8X1^QGE'8ON"M)=N_.,D#3LY>\4DC^9#( 
@4A)T,73-S'&]VNZN=UZW$RGUOC?/-_.T%,?IW]P9P5T 
@]=7R_#M<^%K44)*8YU-V]/A7I_W5QIST@,!3 P,^D^4 
@>'G&8OYK=*W;R03WCY9U%&,-\43C0L36G+0ITPN N]4 
@FS''3"\#TUY(S8MQ;(65A;Z%*]%S;Y&U/F T@4U:M/X 
@SMBY30"!F;DCT'BR$)1:)[[TI?C-B4I'\< ?-H\3'8T 
@K6.[ID*-Y36=%9%%VB^\'A_"-3;_X9NJ[I#L\95RBX< 
@,PSG#'=:<66=MKB0TOU&J#\O]LR,"R[6GL%Y/%.;"C8 
@2PA%MEIJR3BYK[8R3#CN/I!%H%66OZ6<'L3"HJL)2F, 
@U/8)9O:'C5UX_[5Q6$^+)KKH"&<<,6P/3><I\W7W^B\ 
@%XJV>U_IC]D9L,KDB3HT/5GM41G23]!@$(?@U/R$YH( 
@"D_?$8IISB]4''7/ SVFL;JG7ZK>@7FJ[8Z&>PDSS*( 
@ES+%$2I)4AP>461"1^N+!'  WP0?Q4([' B49/;#&MP 
@<T6J-:]UW\<72P2>W O>,R[J8C/CUS7'76OE+:_\K)4 
@8"&VAG$ - M](QJ/T3GE<\7JX/ ,,1)1K5*DTK@X<<\ 
@-D"* 2 $4V5JJ8#@>SF@\[D/%.2+T5S;![*!Z1@C@IT 
@:ELK_M3E)EQG': @GJ#!!-P8O'+IOJ&&*11/$F*<>9H 
@::.-"O_Z3-!?@LTV?';[02'V"\M,W3>C"G?1N9%?RQ( 
@2XWKU?:K@I[:%[-/W>C;E [))9M=UDBYQ4+I%X<@D/8 
@15:T:,G=7TQN1S:%&<\98KZW9E+PD^'^GTX(N9^JE^, 
@' ,>Z@4$X2"= ! 3=DPY[27*4<'*32_%F'.2@.Y",H  
@3+,JGO;'DPE1>W(ZCVRV^<T07?>Q?&D&&GNBCK0D=M  
@0(!GEQ:;,UX)!0-9RJ&B#M1179-P./\WW>\D E4( #( 
@HF!^1&EJ64H=EN%YRVBPLILX2D,U":$4O#0+X/:70<, 
@>W"E)?8RU6OZ(.?O0"$8DO <HK?5^C'L_Q/\-FE3FQL 
@FP^J>XGF-B;O:.HB1>,RAS=,-VLT:"]=[RBRE\0W$!\ 
@ "*#9"G+ $Y^MKD9@Z_W/HB8RQ!4Q;QBX?W#X>56.N8 
@&$[GB+[9A93TY_GBPDLN1[R<90SV1W"*.8^5#)^\>LD 
@5N.()D %6?A"U A76?^$-:F[G_5G\M%"4^2+6:B'&IL 
@":?81*5%DO=%1UZ5HLA/<QVM>G+"S0I%C0HCQ6E![#8 
@(]C9OUQ.UQ)N%W #;;7!,NXF*N4554R_-Q(Z:##'H_P 
@3<C5Z>@9?QB\#H.'8K0!?ZSM16H:$O1D] $EWJ-X8PD 
@RZ^+AANX%/GGXJ<S6]WUGOU4M'1C*J=>B:YCCW2G-3( 
@II,77K#O*W(SZ,A#3_OD1E@ZD:#KX5?POQDBW@8_),< 
@$7R%C+=HJ]<NR>5N5G.SSST)8H;X4!4=6^FH:P^A7%P 
@G2OFM9A< [6NE'R YJ4J% ?LKP<+ :D4'KGAY<TPIY  
@?-?=?"X!W.@:KD:RRX[#*-:2>0N/$A:0K-PE+FU B2@ 
@H*0.2NKM=SM;0^85Q6%7DZ9N9C;O@BD.RXX9Z)R8NK0 
@IL38O;!&D$ ;?<-RU<REE4TGV(AV,0PCO^%-)BR?O[4 
@;]$5MS3 [>A95R!?',=#3H@-L.&/,M_K:J<^L0V/><4 
@%M'-2<54IBR\HYF'=LP&2(%'A?4V=BCN6\B5.(AE+)D 
@AB]SYL=;M5%5G!;C+R!YQT9.S9U*@0W)]DSU8RQKD3( 
@D-\3D),8F=8)JIHF-$TO]I1P./H=>QR!@8\'8YC0.>$ 
@+I;%I_I@J(H-H5"$H7HT15UH!L)OEJJ)_9LRN-)$^AX 
@0C0=/"!YAE8A!N>$!RC)SV%*9BX4_CJ!Z=1#5.V"E]\ 
@7WDUTC2=XR[%*OGFIN>*V5VWST;]CJUPFR;QQCW!JJ  
@'LC_*$'?2ROMMAY#56/C9O243KRHCHF4EY$-P6!&F^0 
@I%M@@;9K*9HF4L':_YE7FRY!M*V!R]=3T2>K\$M+'X\ 
@:=A155<2BH)IMWZ%JNR2J:@$-J:3ECQAXQDZU6D(6#( 
@<*HFCA-*0+*@KU!AL.;E;K]+?L!BI5.7*$WI=+X1&N4 
@0I'B5D,M5X%$T;=R%D8W'I0DT$?>5AFHONS%6*;R =< 
@2?W<XWK[O]4O@:D2&7O=/V*-IR!Q*(+-"N#X2_/O0L8 
@1:&/8V^=#7BZ9$/@.L_K'.[YBS-\!/].:?>CV_KKJ:  
@Q(-8:83FS^@HTDJCY1A5V,)YR/_]]X#BT*/[ C=*,^< 
@SSDZV1I%OV1\I;N:7IHF_&@=6SU3"IV+^9M\ =&*^!  
@P1>X3GF&^63S5T1OGIW=CUKU#2;7Z)?(KC[QR&)G88P 
@='5V0)FRVWBV(FGE'*/X3)A:S^GJ(T1NS O):PF0N54 
@,Y-Z/%M4\D7;U$J7NN>UV\]Y8^L4O-@INI%0Y-G#_X  
@YMQFT](N^COC8L><M+9X%P$8@5"OALXSL</A" ,=(*X 
@L0#^8-LI ^,9,6S"TIH8!!9NO2E;2YE==E%8A?NAC7\ 
@A4QP40K:G$UMQ$-A5/6J;N/5\>4OV<?7X7TQ^RJN!0  
@QUV0_/A]>Z([=X%>A9P=BW =VHD9XL R=L_02F?B9,< 
@HVI#22T/&:WO[<MV;VV?Q\!Y7#V%="R#6U3S[>;6S2D 
@SW>FR?RYUEE.^QB91[&'3IGG5B4\QXDA-G$B\>TTR H 
@4)?MC<\/'D0BUK&O@FPKG$S%)\3&T/2>I35FE1$F]#D 
@0'@Y@$;I@]%_TB%?$7^"U'G$!';A=YA[XX7")2G2(VH 
@O)-4/:Z'-S2J=4OGPBFERK[0>\(W3=2M#SZ<T&,OH/0 
@O[044.)HNZU1L-K3<=!DYPH4(WX8SL -# _J(G/36-  
@[3-9LS\A8#5-X#7@Z@+K'T ('-63X\ RE53*U&UPI:T 
@T#\OMWSUNE3)QAJ<&^,6E;G"AB$0C#:ZX-FN:1C8MR$ 
@7Y0Z![[29/*=M?S'#L(?&&8P:;$"YO/0Q<$=][,!:_X 
@W+T\U1$0L1KY^-2%$?X6'*[ZCV224D>Q?C-TME>>?C< 
@1CW8M2S?(]X'%&DMG2W/XG81\.V W^P5?,T$HTYUNK4 
@AR7D2/ZKIO/I>:U9PNAZ>?$J7XPWH%&CU%][MP:?E]0 
@+\S=.3:6:NU+6\:"RN*$R>Y0)+ZWV=*L@U7-:'. \U( 
@O47T>GPFPP?&V)]=U".KC@W=+Z#V-0H?Y@H[=/JSS6$ 
@YWKV"NDA%!@ ]-A0YT8/9:T=SUFTIE,AO#%=V>-!?"4 
@T(+'+@"%LI.HH4$Z;!+E,F4<S(YZP^$I0@L"NG'+WI( 
@*$YLTRRD62CH*-:/A;ZMA-@*S=Y=T0VFT.PP\0@NJRH 
@P* C+ABT&0D@^ N7/Z@4E00J7T4140[?AJZE(,S&AC( 
@=Q.*L8+"T<21%XG.8/"%0CE%)[BH3U>I9+?J4$S+L)$ 
@-$2TSF <08.]KLW@2?ZF).[3*0^I@Y2!Q 8/N"\/9T@ 
@WU53^(0%9I2>@<!A'7WC?1E13!J;-M/MPK()?W5S9=X 
@2HD5.!K:@7C,"!9VUFNQ)UC\KU \JXOJ1Z-=,QZU4R0 
@U+5^E\;1C$ ,D,QKW6E9W"4&FIN8D8YZV9?E%*@:E5T 
@WNKI/J!17% @\]D-1<"Z7A9Z\,88XPICM28*F(N<@2( 
@N!&H6U1 [?4]%R^OTH!!A5ESRB8H?H 4JXT*>9>@YWT 
@R"24TAL2G++2M0)[I>?4=9?KB7=<!0$W Y:ZTA-B5;@ 
@:A6MM"1H9)-]P]3W[2S24*0-R#E>(,"=DNZ"7Q+"%?, 
@6P*E0EMP7)-56&8J/&E=7G*_)<:D'M9S(@?6YR_9ZTX 
@G]$A]T- 'TU7/7&)5;G%K&Q=>E!ZFF9E!X?P)14+QH, 
@!N)! E:U7BX$J4M#$()GUE7^&MTTA,@&2(@U0$/\[$0 
@8H@M;?A#SG0*&UG24S2BIE7B !5%>!K+4,!"24D-,Z@ 
@\\A1[5O/\[T\D*<J5L@)R<Z>@334)FE"LV%V'R5T8 L 
@5;(_-.TDR#F)7($Q;0&1GT\ [=,#.^6VR,LC"0!S'V( 
@;*X5+Q*O5_X9FA,9572%\+AE\?OMGCC-_J5T<M'A*U$ 
@&N^X1&?2Z08?/1>0N5M1".XUZJ%K'A=Q;>(QNS1I,Q8 
@VM94G9%\S(D7!D&J'??1)_(,(B?>@H)%4Q"?9BW(9NX 
@%DS.?M/LK'Y8)BP@<,GEX4->J\4"A Y!:P3#')6,KQ0 
@VTXA_G/NPNYZKJJZ9H  R/)Q^P Z?2%NHH74>QJ_.)$ 
@LAQ5XI/'&M#WCN\TN6(B3ZT3'1$ /:P+,ZBJ\2?-9]H 
@"N;*:Q]%JK=&@,'K,FHRL&(Z3&Z\"B>XZ-#Z*8V?7*@ 
@6;1%F4=M>%X*"^DZHO5 B!089_0+A-2T6!<5Q@M9>10 
@&W]E%@P:LFQ$>/5%ZR8C**5.81I:%70^EUS&A7,U#$T 
@0!I>$U5E#"<*GGIK?7C96G6T8C.[=2#W2 P#K#!0?W, 
@:,N.2/-SGR)_O0IZ>\=]\!!DC+&S_"3F=QBC_79HL3, 
@.,U(O:2=3M)':^Q417-'[!A8QW2&@%VNSW'AJE)C(J( 
@=YFOG6S/W3NJS8Q/=*PCNDARN+T<RS<2Z>;16HH]%,8 
@,#"^X>B\5#& @L@V\3W2$DD22X=!E/P.R/+U  8?B5\ 
@! !]+MBP[-V!#^GW<Q^C\]JM+^@='KS-:E^N9 M+M4@ 
@SL29T<TB!E8!XB^0+]#;[5'Q+U$!'KA)?-(/)6^+SC$ 
@8_Z\X>0@<AX7X<I'1TL]F$8_TY%"1=7=_2_@8F5+*9L 
@YD*Y:[=;90O2&]JZ@8S?#S)ZK56/KEGDZMW<8VS>E#@ 
@U64(?P'MV*(Z$Y3.4I)WQP7KY=6:B70TK[S%*4,'6T< 
@9BVC?A5+.!+TA817.%X 1S*]'?]8LW*A])Q4HRC_!70 
@'*^4@%_X%2VMNF\9<RW;.$>[U?(VQ>*\M<^?$8GSI&< 
@^WU\@$^S!D[W2EX^E\Y+- \Q/XT@*R]C.E@:RX#DI=H 
@!P .N/P8YG*$#?1OJYR@VAS0PY##BXR' T9^4JWH-F$ 
@V#TC1PLS/%:OF)B*K5LD-4F;R";?Z^;*3STAB7@T[KP 
@'(YY AV 2R0-Q>FK^D- UP?9/D]P5I_D1]K^^F B;@( 
@(\9U("A\%<-0EN619P[DB_6N/%6'C1.X%NLWJ4O-U*4 
@N46\?P#03(!VCDOLW'YT_A#1G.K)**Z(AUPUHFMLZ^P 
@$LHGMVJ>+^7+D7([UM(]/;N+2G[1>*[#B(JA*<=ZK[$ 
@^JI_T(<MU"HI&BR 89[]Z5C<*XA5 0=-U*S6NK:MBHH 
@(K8,;JW?&SP1@Y0&K:#CQ#=2OKY%*6JM,3^D",W0-'0 
@QJE++A<6JN2@S_TG7>J&P'%X.4MKH^SVE),V>G_*A$X 
@R#7WNBD'L^M/.S3BED6K9\NC=OFB ,_.Y5)E!!=MKY< 
@;1_I=WWIPEG'M]^V"@GV2SSPO^TC2-3HUC.^3!@$U)8 
@L;%NO]@9T!U<Z_YJ$K7AW" H7Q=)^K+OL<^;_)%G+-$ 
@>B<7 /IDJ[5*5-FQ66&$R/2/=M,O&A?EZ KPDU8<CG  
@!!(3-S(@[J# U=EVJ%6K;@[W3"#D)PCRNOXE2PWT(Y8 
@+QXH7N=+B;(P5]QJUVZ_#2E$\>TM_B=\8R %Y0,R'C$ 
@B?21AT]Q<FL6NHE.1YG&\ZX;:FDQY"J>ZNK -H!8N@D 
@2;-?\_21PFIKZB<E)=0\'ZT@E^:W_<&47%8(1(WAR<D 
@/#PEY3K*HJV\ZQ-Q[0S?#;Y\Q[O0:< BF#;!,-[FOJ  
@N/IP2?15VQJ[5D3Z,AA6&LE_FU'' +PKYB8W5X;3VQX 
@+M=+.N>B]4DVN!SF"<N4P'FJ\HX_1H #:;E?LPG=5[4 
@GOPG-OWE^?VI%'MJ\4W?17Z3 R"#QNO$Z8&JUHKMTS< 
@AT>=ENZ_$\H=#JIW>8[]8:Y374?]5G&:QU]O95P"3YT 
@LH#YUBX'*629#*NE].SC4=V%YH?X-0:$Z08)&%J<U68 
@6421*,Q \Y])PFF"Z^S2;ZR_X8B?$.!?.?GFC:F+@/T 
@;>9%2;(TB:(8-:-,>E:D5WB1X%?B*)QC".4'4DVU(N@ 
@"Z[.ED85*U*+,L.XLZJ1XES3V['(AJ=I]3!L0K=4N?, 
@[1:FP(>2X#<6GI,F&*?&/YX_EC#@"OW#810EI=!]6F( 
@[X/$@M^\SWIA)'YXVBG90-@P00L81(IG'0(IBHIA2#  
@S11 *[=S7*9@K[&S"E$RC71NY_X7RTD/*3KX$3O[HR8 
@;L]+CJ*/>;B]UW#__^7G;)KQ=(_"AAH(^@(+YUU1$'L 
@.#.(=82H5:?G"/5.9[CH%LC-)V_JI85P ZM02:5]474 
@,?&]LYW@0*G*%WM?3P0T#*2!([QAVK9P)10\;&*74H< 
@]\%14CE+OF'^%=0,.X9\ALOW[R:**X_&7P_+>D*\:5P 
@4$)8++V;8>LPY%O-3BHI]A9_7#YK-?@!NM*1SXN1-04 
@X[-]MZ[NJ6CM0-J2,>XUW3:HM/ET(LL\?6&F)CL20HD 
@3CP$E@;)6N BJ*,L!N8-'E.T<,C:L3,"^2AC.U4G+J, 
@9W>X/ A*M. 9J( 48\6_24,)P!00-+$];G(>8AWZ<[8 
@91 N;9+5@/]0RL7D('GV&Q^LM2@W$ J,T,:JQ'D?)K$ 
@U;E-(=+)ET*!$^3:ZZ+_%55-+%18)O0I$0T+!^N-[(0 
@ /#"5H8 @_2P5":):[RV(@XL@1>PMED]FF1-,D1H->( 
@3.54D%+")KQUYLNJJ!X1N8.Y,(N 9ZCJ@6NV!)[_5?D 
@>"TE#PB8.STS7M+M@8D9Q\ZRT9JG(SH9T;[@]NQ4M[P 
@W=2[Z6(Z;?DEOPJ8(H\H@CGD*+RM3;7'BTC;5)5_H", 
@8ZO#"?WD6LQ%,HF!3-OMNX-:=J  VNT(HD@*.8U^]OH 
@L;QETT"N&!$'3O6U_7/FHT0CSAZ)::[C=66J,?!RJP4 
@7EUR$FIN*;$Y&37RTN>Z]0-CTFY]=?)=#==-P7\6*@P 
@4!J*>7\CYVZ[BF!2-+2TK.O+#!6JR)EY4)9C+21K4VL 
@$UBC(>/_9?B#>$I:M2!G=F@2YJR*<OM]K['B91Y:N0H 
@4VQ=D'9E8W!E7AP8VL*1? EI8L0Y&$-%FF43>4L-SSL 
@;D]M1#:_-ZW*T9@0L:">[X^E@-X0VLH]8EI K.)YQ08 
@C7TODVJ@^N1I^>JV8<Q]=&F;SV[2$BS(.F:B 92B2+@ 
@YV\L?TL7DF,3/)'!A#G]PS]Q=4$KJ-]0?!\,D<;:;;D 
@T"6-'(%:83&<?]D11>Q<C=CE()KD:.#2I[V8N ]/N<T 
@W:Q:_!Q.C;"9E2_5+PX<9E*C YW"!*>LSD.F3P-'Q"@ 
@N,><;T&[>"^G>#L?*^Z>J.W$>/CRC%+.Y$B+$RG^3TT 
@\-<:ES'6Q[R=*N:^IK>%6[+!FO:')?H$T6B^PWD^4=P 
@M5_XT[/=9$ZLZVJ;GVT]P*O8A*%U\*%559RC7 BL+LP 
@UE%3]S8PVV&CMWB/!S=.>!$9BWJ/7 ;PTO1M0RP9LF< 
@7#4J\@)XMFTAADWWRS:H&261(@DI*%*O 72EET'\F?$ 
@IA0[-=^NY(/W%5I(5OR A0?<M)3%-/0A?_1W%-0J:EH 
@3%"6;$Z6L6I5C4"3-^%IGH#WR<V!P=-*DA51T,.S]:P 
@PO"F^:6*GR7\D.^9,^D>_@#>FXY3LD?"RQ(,9T8D9I@ 
@D^N^DJZH%VB)]XH2G7X5,XCJ&+*75$IG[U&_WQMET(( 
@!!D1S$+,-(4%64*:8K&D@@?JG.6%8CO.;RC<RX")+/( 
@$TL)3OAEXVL-E6Y4E#FV;'[Y^<V@'(;]C#T=DC%F&%\ 
@)6[Z^W8?CB <<Q?,@"JPDZ"E+D-XS-#NV"<D=+&] NX 
@,O@)KA;6B3:K^-S<#)XJ2H9<<>-^#GD?D N#O2C'/2$ 
@SU#4)[7]SH!_0\!_GB<',\\< O?I!C4QA2#*LC[\;J< 
@BL,%JK)\'.C&KIK[#;$FLFBX:IT='QJ,(HM<51E66(L 
@WI]P8=Y_RRQM]D#!5>I+'%"J/'HFAZDPAA5FI3 -H]  
@7SQEP<VI##KOP:*6;Z!Q>,G9]"4B$PAX]OA=D&L>9DP 
@]NEO1.DNF^E=2\(.3MECEP1-K/Y(WD>]0I^8&&TJ+ZH 
@7!/<FJ:/>S CN+:6%H0A40.9*UU$O*MA=ZZ(*6(\85T 
@\0AV3WO-K>D@V/U'":U; J5\;[]_M\!XI:3WW]]FE_\ 
@H"$\OPF[ZF&D%KD8K4- ,#:#-PE0+A!<MZF+J-W;B7D 
@!(BE+6H*_1CS3E$@&)5KUSLZCA]!,V8;NEX J,>0*X4 
@]/G?RX\7\.=Z4E2=NU8K_!GR!O?D2P1!6 @N&@Q2NK( 
@R"?;8YT$!I8U>WH&( "()ZD:[?4;%B256*^? @O0$V$ 
@\CG1)D;]4ZQGGF\17<@_J](E*Q8UP[,DE)+%***0P_L 
@0-$FKA/-.C.$4R=+95D/ZLQQLW[^%5O9NY*F9A/>1E8 
@V7W%,\Q.\H,[VJB3'%T*XBV?O577IA0DIL)]H>C:KTH 
@5#0,%D 4T#JMN#W)(!E;':JKZ1+.S0DW62)E-P?IU.L 
@?V>$&G[^B.%O5'N[A.YNYV!0=%#6D.9=N8R2)?[O L, 
@-H5 (16T.L:L-;/4VKKA[/MD 9P\SUM#9 QYR-5-,G4 
@'?M1FI6[>E6I!-Q@"Y8@;P_PN]<%D5/SVB05[/?  #T 
@P!6 WN ;$6E)%T*##6"OTHMC0;L[ ZCH^(1;;Q["T_\ 
@M85Y0%QH@IW)KA4Y=^C/J0V-Z&)"A=ESHST[G7QM?%8 
@\)EGD)_O!BS_F2P0)<JP!KO4!N+(W8T%[7""P6+Z2)0 
@+:TG]X1XGQM*7F)]HTHKT=H07IRS@[#.59RL!J'WISD 
@6">L0#()R-Z=/'4JT'* 5LM&*DK0GN)8K.W>?4;GONP 
@31OA'>J$&1Q7EQT8O.<L"I21QCCAT#DCF,8L]E-A?ZP 
@QI\VWU.8*?40*!;4:]@^^'&DH-A-W9S)))1#<6ZI3 X 
@-J8^H!0QQU_QP&R6[D3CKI%JS347WL/3+T)]U:\FEV, 
@)LG+.L5%/CY""@N^T&+QTN-M42O\.0Q<*Q#Q;9MS@08 
@9!U==97^"^*A*$/H#@W*2W>!&5Q&\/G+#44;8!BX*:( 
@& 1&L@Y.?+&_?'6C@9"II-\Y#[AGII=>=?UL)T?R[UD 
@WV/6/98B*K#9-0*<^6BU.. X,>P@ W4N7FRT2\RU8ZH 
@ELD:$G'.H".^TS8Q#@SUZ7;$"-<5;?N+ ,^(T2P%]]4 
@.<W!VQ/@"Y=H"R"E7MIE9W0^T>\T-MS0VQJ/TJU?A@T 
@_6VK^\M#&@&RL48#F=4P6$@&4XVZY'*,4KJ74CE9./0 
@,>83(?Y?M 9(EB]A6"\S-%K>*7UJSZHQ-8.KR_#T(3L 
@<>55O_"<+C_[=D,54&J:O;-WM1"3S]PRC-P16+.RH4@ 
@RPT@U&Y@*&SK(84;=53RJYB&01C#0:'P*PU"P1+Z2;P 
@,':QB@'DGZ^"ZQ4_XH-<3\UZ';\H]=R+DV'*$0,7$!H 
@^_*^P.46L5<LIR"&@2*$Y1H\@4;(@A4X4YWW[*%53$$ 
@BF>(?]1'9$;9BY<-2K%\*J! ?O?)Q\O[MHFD>>_S62< 
@4Z&V-%7%E9:- !%^0OJE;G.R7-?Z-XZW5XT4>,3-B*< 
@[I/'#^(J>_(X7\K83&2ME?ECHF1)OW&JF$XA SYH))P 
@J5%"&:U8&^<=3?,X?1(:^?YVH5GK0YY7;K@=&%XH>(\ 
@*VX(RR0S*#][9I!:,H Q@(*UWE5\42 U1R>:'./Y>G8 
@..Q#2W" *RZU@R/1,U_ UGK&S3$<G1]</^B4D21!,V0 
@)\Z<E*P_X@3S7B+<&9:C4N"%N'_V.\))DP15/_KP(A, 
@6'N0&>2F+!-E+UH0QO</V4PNN*;-Q*DCGQ<".HPJV X 
@I2&$^;E%NA#XO9"_S!4,!G\5?C??(XE)[;K7^,O5H38 
@J'-C>S6P<QWB[J470$5BN'\'!YVW ZU]:UAY3S#-V>\ 
@3HNYN%DB+NR9\8=)3:8>60MCSJ0_=@@F7;L>7">&>\8 
@=+H0@/2NE:DZ*27+4'HZF>D;\&B2_QTL4@UKXFV$&Z\ 
@25@0K7*RZ"V5'A7$)B!7BL!99CN!?1&+481<7!%F &\ 
@3&LY69GK$]OU=Q4[UWCZ-;.T5TFYH<4ZE"SRS>2$@^, 
@%V'S#5A_2L7/^MA57XX.[<1CZ!>;G-N^W[C)>K#DQO$ 
@X5RXK4+T\"?I_XDK@97NREN7MZ^Y/07&P47!==B8P54 
@E _5Q])O\",F69)^XQ1YP(.ZH.W'"Y8MBJ=%,.%LE8  
@3>WZ]\%B!#,1"8I,@7AP"#NN6?R4_$^LIBCI6#G]R\( 
@Z[</#^$^ AO*1?4!GDQ<U[ZJ!JO3@:<ZDQ[18,C=M1T 
@A<VHA@' IMHZ%[-.A!!4A%I0LYN+R7'/866B1\[7YF, 
@]PYJ$VN34AE)8# >9O_$RRBJ@7=3  /V1$_Y(<X -5@ 
@QY1C% /_ J_>Y/"P'?^236YTYS@@I*3%O7G1[85B':P 
@*)R]\\=T#JF&TN"/JY[XQB.#XI7 ?F"M2T,I@'^#, X 
@P!H^W],&KWSP5BIZ"55J]&=\LIC6^3%B,GF5:;.>!>H 
@>O/9TV:5$5TRA4;4?9A!_XXAW;@(.)[)]X*OB>F3.RH 
@2+W%\#Z(P U= 1:]X6YB[("6E[%PA[X Z>1OU#/!?ZH 
@I>K,#QG#/6S_>$DJT[!0]\UU='&W[;#TAC?P>"3:B-( 
@7UE'Q@C"_T)Z);RB0P;H'--&:+D@"4Q!"H!?5SLV3.4 
@^VA]5:PP(AAI_C! #,;DY/@68ZFA450'97REN%52/O@ 
@JPL_6[$8EB!J\\Q&!%H4\WX83YPI7KMGOA+J-& U_B\ 
@_:(.;&$X;#]?>";F@%HPO &<<\+4HI1-AQ:HAJ@Q=KH 
@Y::JX>S4FX6WR\ZZ6TKCHVVX!;^OGK 0X:W(A9R9&R  
@NY5RMPVZ+L3:-#66(1O<'DH%---<DL)Z \!G13!%(O, 
@#O*$:_9%FU_Q_G2-"DFO,T!0 R'G='0%@ 9O[P.]JKT 
@55<+/NJ'6]55Q # 5[6G4;4'[S#_-!!?0]D)G4M=Y-4 
@@J@0*H*VHUO_T315!(F/0?>>"=_[,+XN+YAUC]];QXL 
@DD&W:8+_Q61K^8*Y"'>;L7_FAD]SC@CBM%/?]:;"]NX 
@V>1WM08SD7<(QR!U:7*6T9<>4A)!.8.WX2N4'*!9_HD 
@K/P5:WT7? [OXZW)M[A+;%+_4/>[@3:D-D\@1)N#_CL 
@(*9BPV?I(QMY"%)YA^3Y]U?Y]?JA*KUL"_S<>=V[C]$ 
@78!O"R0E+@K<F.I$^Y4O95H@"I9&W;E<8(Y^C1=BZ&L 
@:]$31Z!) FCXFP@=IX1K5KD-7<67TKX6E&_&.-<PB5\ 
@#M4?%AO[I^FG[,8'#%?@D]<AOBWPO.O2+:$IX-]97^L 
@(+S<*HV> #3."U<\-:KO5WC08F(<AO"8,A+5QZ$C_6D 
@O]\M7/'NE'' 40<J2GR:#9HJ5!,BEP;B]&VIQA4.J', 
@P676V\G?)79A?)1=PHC54BR>/;$;,?%G0P&ZL/SXDL@ 
@2ZP1,]J2A,+  GJ-CN6A3T,- ]HN.RDA<$Z,6?CU+0$ 
@$+T]*K.&LVW844#-Y58=(&=,\1G4]WR QMG;7:T(Q:H 
@HG2,6@#K>(TR^L-JLX:8AHUWO2I@69EP=Y6YVNBMI(P 
@_H>\GL@Q&32NY?B'URMN[;K<(D\[0[4T)ZN+7! +]E< 
@)!WM$I9 554[=6)+D*DU>H!7]Q351MHU2LU./CS?/#H 
@;(AY*]JB*N0AN+BKAQ= 0U2+ Y:5?#.>O(XE%K(M*R0 
@1#"X53L3ZML58-YA^,/=76OV"OKF!D[DH*R!!TE9)+T 
@ ^+Z4$3S@O?^40'4UC1VDL"H#16U+RG84JIEG&.H[OD 
@0U^/E[K)SM$W,-,N.1B8.6 ($<S])%TLCG4V1%[88ET 
@2=VW^&L]9\7RN<%7N=3IEWG'\"Y-6J(;BXOG\Y=GH[X 
@3EP;;EF'$"HJ>1:A0F\0R^ .D>\]QFX@S!$,LO"@='H 
@Q;LG-*:V6W'HM,3/_(0W-7E#;R./M&5"'J2!W#.?RIH 
@V%I+(-7,A\A.+7^CVE2_<.9Z_D[3HFR02:HF]HM"T4< 
@N&,,=/@+@2"(ILQ*^E0K.!#][C,#!U0<FFCF:+@#UA4 
@83IV[!K^X3:+W' LG)Q@HT(^CG;@8RN%W CF'@4?!$0 
@UB,"XBT[Q.6DU/C3<;_A&'U).E6&!7'^^I80-,12L.H 
@A,9YLC4QMQ:/[/-ZLGIL3&H@8M\&M$YHG:.QFEFE8D$ 
@I=1^[DWVES/FM]SD$=A1-ODQ&XU^2P-,1;Z^KP\+?+H 
@)4L;Y\:*D7[[W5)0PJ2[)'P $8?6P<B9^842)E.FIND 
@_"3L\1FZK;6.GZ @^I)Z*%:@'1OV*[ 1AZ):((T+IP( 
@26,PKXZJ 3),V>C\M)<I4Y*$?(B4[([]]+E&H6ZP49H 
@[UW3CH\L*F;> MZ#;RI_DEE.%39B(CUL=O4IK)S7!%\ 
@R=-]?'MGEN"6R<U07G)G'F-26&&'#C8H[8[DW[N;H 8 
@-!):N/T26VH0/D_L4S'%/RK%UK9U=^;3B!/6-/@^TA< 
@1%*SBT*11#='\#AZEG3)./D*%6]R_2&E?N=\)RA]^@T 
@36I!A-[)-M 7T^A@O"7#81A^\P=H=Z.YU1Y$@T9F&.D 
@Q;6#AI+$K#S/147KY+_ZV6S9ZQ+![/#ONPUE[OYPUM\ 
@H5P+RW ,KUC2)53$!)=&@5:A57SN>RNZB."'VB]P2;< 
@H*J7#/E\><1L^"/YV\M2.91=H\H3@^I^R07,U5Z!> L 
@" G&NM.%L9EQQ37"/KI),$,EX9H84?*G*Q(Y)'I88RD 
@0Z&F"=6#H<THEGJ/+0S_5A?.%@PL?!LY"1J+C\&PH(P 
@%8[C%?B2&46XU9:0"-B\VN,4GE12LUV_?$47IV*'FC0 
@6V0.INT?JHI40'+5UJ(]YPEX%F5E^4I8R0A9]F[FD6P 
@^@=>!%N.6&L@KT]4635#'1%Q83\3_IG,D,A):91_7ZL 
@M^I>!22O4 JNY(.8K\:S#NJJ54EG-%N-_T],0,?N*]8 
@3W<X&DQ0H='Q]87U],ZKW=&"S:HM"*ZUTC!PE"N7GKL 
@,\7D3^ $CKMG0-TK.YBSL-O<+D%PPG^</5[I8LME+=@ 
@"17)]8MD,['Y.F*=P'J]3.2!'6XPOX^=UV-DV1EEBA4 
@F?1WL*Q'^=&Y\EG+B;6LF^L$_A"$I[_[$GB'93(4XTX 
@Y3X19$'?\1!D-P(0*T5^.<PKM2U&@E(7$]J3S#FQ!4@ 
@\G&P$'@+><F:7].]S0CZ-77>/S)_\2^?<=AZ<^&R&;4 
@*@VC$4AN5A+?$.JI8-2W[6*3"(>12=&)I![C/$*[R@T 
@+8E;0I16-RR%XUG=''./$Q_+@$UACCXTN[C&BL*J'J0 
@I'[-H=F32=$V!N> BW*46W 2[*N:CAHPBUO@+_8PR5  
@@YS+%8^O<D"D4 \]\/SN6U!5MQTOX"/X7#NRAN(*[-D 
@NG@P;V<%:#-%J?LU(;^LB D,TP2RV#=_.=Y31&R^>%, 
@WY>!EU$/LI,YFJL_H:E5Y=8)^M@H-HV[$,88/P^*J%$ 
@Y=L)4.KY967YV\,9.%A2EV2JN!FA7-BE"?==*]CPQQH 
@)(5GO_L4>PQFU#-Z/AA3!"\ Q@W=S$L %G,NFH0(7J, 
@4$81DG,G]0TI&J-H1ALW2V#!89Y>)W(L:'B%;))B8TP 
@%I /Y8_OY22@EVIL"CPDQB(W[7?L&P#EEM'!*S6A]GH 
@/FD_"Q]. 5&-4A;;$:Y(WR/)52M>T)J,U)"15IR8(N  
@U__[H1"9V+)PNE$&?#!=_R:=S, &'IVFL;*;\<L2#R( 
@\4G^,1$]-%%XR8B13I@U] W"B91N,.5*T!!@_C<X12( 
@3A[=YH2"%G<Y'W;TMXW3&9M>+.:G/JJJLW"EF\120[D 
@[4,UVG7-B[!O#);-5'QB,%;RMQ92#01\RP>60 %>WR0 
@85A.(ZBA^2:1((4,X[OQ_:K5\#W?1DAD4GJ;'@S)+S< 
@/!_RGAWM_@3;DY(9'*,WQH7,7G/<#?R#.-HK)/8/-N@ 
@V^XI,%57=B!80PDN>SG>2F8JU^QS]8# QSK8$QQIMCP 
@"L)Y].VO=6("T+I48.T.[@$/>P/P[V0OA%XV4M\UKK@ 
@%,3BD]4@)L!)=;E5MV73V5V\8H<OT'2FV2&8N@^0BIX 
@45\WVJ/*%XM-%$RPK:JQLC!NO!S2//H4BE6U3\:MTE( 
@WNO^NFB:0FX)^)_2'%B-48UL5>OZ/,>,5.3T+WMK5X$ 
@,X!W0N\\UT<(JRZ8=]N1ID1?LSX5=.G,F(TESVOL@_L 
@#1.O\AWF/4C' $[D:_2U6=^K[]=Q=W/@"GC[G[NE3X, 
@)_/4K'E7^B)$&RR,\LM)87@LQ)OC"7T@\UT4G+#@4@H 
@5WPN%^+^0WF[3S_V0\/"AHNE2;63A;4&TANOY;,W@U( 
@%5I-+BBI-;"W2B>E3$,59@$*-L&>/ E7J3W":9.7C., 
@Y8V/VJ.:"E$WDXGSN!-IEQHG!',CQ@H@F]/AH"TVR<L 
@LF*,,6A$D2 "4TEY^5QY8B,=ZO'AM1I%:0*?$5:U1.( 
@1Y6D9^B7%WM"9J6J3X@%'O74IGHE-\0+R4]#*$">SN, 
@J6FEW%^)YF3Y>>8M&Q"F::"2HB_H0!JB)9B<)T$2+N  
@?DG?:BX7I\-8;8<UD;KH@O@*M=_V4YZ.G%'H[F&8NR( 
@!/P\77N<Y-%* CON)_6_2'_07XZU:^A"GC%#7'(O6O\ 
@"'"]/BRG&N?#L.$4N8FY21M_N54$1Y;,F8 OIB><F\L 
@D)SZT3?\5,G:M34;W)P_JU8:W:L1*DGL50Y8*OK0)SP 
@^>TI7-DN<HC/"2W\,)>V.S+Y$!&H[(6- ;:6(&=FP1D 
@Q[*HM! 4]3=%#88$5XV,;TK(*/8*HE"M^Y3FC<KC*C4 
@!@%AP_D[!LK(!9 60>CLNX2-9NU2B?>@Y?*#-/L!UU( 
@X8Y,[S#/);V!@6P&MT[;M5SV+B-\@PD/]9?T9BCHDE8 
@W\YRMT2BG>)"RN30W+)#[OQWZS3V8B-L7-VU<9I@AL, 
@T(PVD.@9=LSPW#]>+G='<-=7B ^,'"^%^GQ0OK28ZC, 
@Y?0H/IL[6WJG7Q(Q//CS(70"ODT  /?]Y<O2\8(UFG0 
@6>%L7I7"\+&51%&P#J_"B(/?G$J;\<")J@_1%) 4K>H 
@5,;,#Q^'004Y_@2*K8D'#5*25PL()FJD,F['8Q,?/NL 
@ 9&499F?$6$ S#T8ALQYX%"O@MXEHI..FH8\KHG-%?\ 
@@'ZX"6MHK"HH-7=&E*-KS"9=FQZHB$9(6KW4=\Z6^A4 
@3VM<8#8.WC)=E&L9& \4G*_SYG&TO@I.GJD 2D 8QHP 
@&!T_K[(GA9ZL6[S%5VFS/@00TX49GL2]UW<HD<[Y:YD 
@9CX#+".-021^7$*^:BU]T16%")W"WHU2%C8F_^[BU^, 
@N>R% '>!",/P=Y\/N51I &*1.ZNVI&?FN8+H^/_^O74 
@:[(53'!)Q;NX&N@J))0';U[GX\U=R0 :L/L=6OXO4.L 
@O/AJ9\N%:_"Q0@C=,ESH>Z=+@LY \V6HMK!FR%#BVA$ 
@(9\4\8^!?= _L=[B1*3?GO?]W 3DP-I^Z>)5,QS\:^4 
@2DR!P:8Z$]O5E(&S4DF"64#>]OGE<G/KS>++L8;9IAP 
@(7M)'EMI'58)B%I&3+W'$I]&V+:< PC;F?8"%I_-F\4 
@&79&/4T$9-AMH6CIK"C)AQW>:1[GUE":X0)8,-W"<RP 
@&5X$*F6_>8:"IAFNW)\ Q((MTF/Y^<(H$NZ#MG8R<KX 
@#4\)BW+<=: [^OH;DINY!+=19=BDYRB956R$D8HX<T8 
@<Y;5Y3K,59\D0K:IB;/P^%(&*LW:)%-ZOVCZNOY1Y+L 
@X[1]<3[7!-PAL)*](WE.L97!1V,?W'99*&_7QP[/[LD 
@=I@>LZ 5'']EJYV>!B(,@4&*S3"3N'4<*H%"8OI+O'P 
@\ [K>ZX77@;G7Q_7H^(N#T@JV[]/;SM:J>7IY<=H-MD 
@[F<NX<9=8:55NQPRU-_53,3>/B(Y:U5@;[U\SQ3>)&  
@:+X] 23:X!R9(MK%Z,9<0$&+ZJ;-481D;YCW)84=:^$ 
@;KG*4KI#VBCXWZ%R/*]0FO6*Q4J<#J_0VY $#T7V39T 
@B'%DBP^&T@FPCF:A XW*BL\<XU$:1K59@?%9TG,VW P 
@$UC5MQ2&7,IS+1AMW-Q7N==B<>>.:=A5N9>"T^_NT<T 
@=C"^#^X7,(QWRII,O**<D%9T[)<*!CG;BN>]T"Q\55P 
@)O#G]((5%@H*^K.'D<G<<Y<5 0GBXADBQ*\2)=PW5/0 
@\/\B5Q!:N[B+N]ZFK#&VH4SQ$R"]%F[ DAG-0137:FD 
@(@*W++@QJPH=,RT-9J=8IQJ&I8#]]/92X'E3+T#+QJX 
@XW*?;^C5PL-QU#8%B5G,XYL5EE_7_=%*MW :*&9ID>, 
@EK)*'*B2X'4WST)V\GR5K9#-V,LT<J =4*,F]MH+FXX 
@^>IW='AS +1 =?'4_!X"QAK^%9+-K,PC@X]LK*#!L-4 
@-8/_1);<XY>;9"7H#.#.@#[NCW)1(;G9M97\3W W5H( 
@Q7H@]OE6?Q9!%\'>W1VIG.,D0FT=!LY26ATZ2[K60?0 
@,@3SF;5.\0@K'2 GD^.XU= M0#;(&:126 F^_O/4F%@ 
@(U+Y3BGW$'8%R<T%IR)&K EBF.DE!$>)G(]%[G'>9*8 
@G>,&60\UUU*@$E ? APY\!Y]*@8SNRH3E/*#@CVJ8/@ 
@/VN2!6^! 3UH+$K8&I[G[/9$?]?MD2U&N@<5:VBFI9  
@!(2D_%<09N3)GJ3;ME?6M"X/%:7@99@!&5UUN25'\?X 
@TJFCO.K-OP,#G/T[*<%;K)"L2=0#U!BWU"9D9]#$ T  
@C$-H_H[WP.>139*(3ER05I055!#^S)'+ %Q*(&\Q!/@ 
@:ZBGZ\KS)3(2?[;Y"OU)&W+?T@MGN" 9>C3 B\'MU(L 
@@DI :6,/;HX"H/2II/4$D"94I=>'+V9J.(O^$>>;V7T 
@421![$PJL-L+K[;(_>9];\ >$6?4<_ N+OPC#PF6R?L 
@$5JM[7TX6?-2(&UI>):DUB48]'S(Z.!GV_[&;@C_ >H 
@'._[_!:=OCZ.S[D^HD!"N%Y/PWCZ57BY<GY4'"4*<J$ 
@[UH@,724_J LJ9*:TML55+1\'8L.:#EZ9_E*"]J)U-\ 
@2-W%KJH: 1.0<*KG=6!$.@L_G*Z-RDRN*W_P-7GT/)4 
@]_F,Y"0#9S5%N];#*_W@^A%FG%/DZ0<6"3;HXP8OF8( 
@0+,<KEU'H&O*_ENIVT!/6O0-SJ"\C]AB3"FT)5<Q8(X 
@-W&'@3CA)+6(94<S.ZH7G0O!J<A:7<$6WEGUM4*QT%, 
@-L'R/KPY!):N9"E+.=<"\$4O4=MA[JBS=N_.XNJRVFP 
@3!+[[(ENX3"+)"0OX[X8^<P0$UJ'>63B@%1DE9I=CLT 
@D;G/,=7\H"@_/[!((C*R5Y*K0IMH%*-P7'G\2SMQV/L 
@6S 6*+G/.<0Q9?D29D[->]<2YN555NTSNOA;/2BK;MT 
@)L"(O]YQ E? ?/^]!G<^44X'M:_L:',_M>;Q/DLK&$H 
@95UJ^7HC*<6.A>)MC_:_<X]B6R?.A(;S<NXUN:><0;@ 
@7C:);KJZ"&7'?RV6"F!#[667(9'V^\3:ARBKB=+&^*L 
@: L\' ^U6@\;#9EUC(6\L,H?6PSJG+:9%#%D_@WZ(7  
@6ICV0]<#ZYO;<]W;L?9DC18X#>-)Z/L2^(2-''A>63@ 
@([_%.-8,=$<\!WSGUMPFAAT?*^]4US#\U:XS RW2# T 
@%SM71CHS?:T^%[S,/6!(KW@!9WJ^8URS$3^: 116M=( 
@;#B$TXG,33.KG+T]HC<#&2RV)^"]HP-)*%QR!U.]&4T 
@ N!3 ($#><,N^CQ[2DVM6>!8VR,_XT5D<2%NX\]O%3\ 
@K]HCVQYE>)9/KT=@$O[+0#"D/"1.O!D=)Y?N'!X&#E\ 
@9S&#>!&Q?38=]7NO%T!DY9GX5#?6@C7MZOK7MGQ)S0T 
@,[:X4L=7D3-VY_CD@(VWFK&RV@K]-AL7E6QRYP+#158 
@RV'/88$H,)"B@ <\A5/M_T>G*AZ#-#!N[ $K>>,L^*H 
@EB,;(O=.?2E]"Z>\H"X+:I[_@KXN[=2;IVB>;QUDU)D 
@!)>YLMPK90M!_$999P])^D=[BA3@:F6)EER=$E;>\80 
@'I1A(:0TZQ%LIZ#!#I!7<*H-1^KV[V+M6F3!OYR0KR@ 
@],"&P<(8$4"%8R@[U1H=/6MZ9E. OGYA1&,-EE ?C7D 
@"6O,].\4&=W!3".HD76Y!?L$*A*I4^ORTQ_PE?QH</  
@%Y_P<(Y._-U6^"9.5N]QGE5=TSFR3DT0C2^:'%S?0B( 
@ZJE;&9G9W#MKS0O!V!^@NJ0NAS-PQ2@6PZ4K<@36G@@ 
@9$[2\_A/&_*-?N2- Y-3@'O:^*K8-KRBM3/G.QR\B]< 
@6XHHTCQ>;GB,W94N_M70T@J:XGQGU?,G)8-$TZ'W+/@ 
@6L..KFH?+E.V6&R!Z4M#^!\HK]GP1QS@.$IN<'"D+NX 
@SFNDV7W:_SHI&#$8$5!W7!4IUWOJ\1QY(0^^[E=DSE0 
@"]KM;1/1&A23<AM@*DE#W0$P<FE2E?[OI!%?NKHEYOL 
@=:!B(X (WU/RPV:S)DGOG.UD:-O:T!_]AZ(4)/';-P0 
@B*G-2& BIDV&&EL2CERZVF=R*!6FT Q%3F6!0U 6"C$ 
@,"&^CW$%:TF<K\_Z?;N,XP&]RT1YD.C"#]<+0'ST,G  
@TSZRV.9K'YV_?T-);;!V]Q'BRIJRD#6@5W%[/3CY[<0 
@0/#[3%QY[TBGIS&8!ZY8T9V-9.>AB+7>/C!;-:(@)Q8 
@ORPAPD'P%XNAL\8 T=26+'4FJZRJOB8R)LVG0VB&C*( 
@!8 N@.<H$.FK^9;G@X/5A;,:J@6Q=GL_K+A1H,D3$'< 
@4.P5_4(E3#!F]CH/XIHMX>/889AGH3P@S^X59J6<=O, 
@P(I#F]PNA=1J*]33OCYSCS0.5M\9N$H-3^W.AZILW64 
@[^"]S6OD*VH_< U# D%^6&H4,FD/!%JU.0V]TR:8*ZD 
@;G6?:)T]V (1!DJ3E_*%8T>$*# 8>6X*TZY</#$T\_< 
@?;?X]!B]/YQ*!U,,$B1QG.O24LTFI'/?3ED%BQ=7QN\ 
@S#-["!F+F6D^/=A1@Y15AW_HWO"K.\.8&!/!/FW=DZ( 
@F.^:3'5KOSY0R@!'W,!+>&F8\HC4N,/:SNZE#YY\!50 
@<5(1SD8#8?%["6!!'"' ZGE.P% NE&V^?T0/8KT^=VD 
@Z:SEKACNWSS$-C)ZV;FD2Q%,2!RB<QBL3_2?Z.%T8K< 
@HW'$;TCDJ&X?R@\K=Q+*+2)'9Z@JQGRQA)L3%[P:6D$ 
@DHY8(;:.EJ5[Z!]]'46[1E7FZ@*HF(;CNW>'1]IXG30 
@TNPFQKW72%EL75K$N12*MF_K@6<B96%R ?L70PO3-:, 
@# <>G]B"!_KF+D[O20_2'XB#5U(3S<2Y#IN_)_O9Q;4 
@6R(MTU/NK!W6S0RNMY+)4_0*FPUJI@B*5Z78>L"BK?  
@H1*&TH.ZFT6+L*8C.B@+$<.62$9$AMLX>@E?5[,]6"4 
@R$/5(Z[2S"#IA(6<F^J,Z-]RT[CJD<-=[SVB-!IE_:8 
@S_<@PP+W518):+"AEWJ@N>_-O(S\#PH%K<Z9YAOUG"H 
@OWYT[&/DL-!.1WB N:2"-RMN8A;"P"_VN*A-.W$/IT< 
@HR?JJ,Q!AVHI*301"4K\-$<G_.KU S8:OUR3":Y+%*( 
@%<0,Y9(IE]J]J4ALC\:LI#;B756"3O1RT<_FX)PT7G$ 
@ <<RFX7E'-B0-1!]^]:ASEH8T#Z;):@?'O"$VOF#@KT 
@?M^"R<,#GR.P6,/C_]4IP&+X'MN&U%%W2=&A0XR$;\0 
@:CU<_&!C8>:0D/R#O"!2R$E1#W9@;W9QA:"?MXK!9'0 
@1-HBN[]&J>"!\LA3&KJ7$6[",U2:$5"RC'\-^,'C&G( 
@!5/I48%'GT<X*+\%#%/0PS4*\\1[=.V6#Q@@1TQ-A/( 
@O=11OAZM6]B0<B8E$($ZTG[."?DA@/OW39/:6%#.BX  
@3")&>*:/=>J,: !-7DY!+OO03E;HHXUWK\K6=29 <'4 
@!WN36G+C[8(,.#1EO\]9H@A [@AV5U?TI:C*WDE=<#( 
@W"17?5:MKY4#MPX@:*6FU_)%Q)J54.Q]&EMJS0M&.Y< 
@ K^)"O;5GFP0A_!4R-R_"L*S:CZC<X,<)Y))O_S+XZ  
@Y](XO] YZ*#T6PD8#1'<F="PE/:IKCU*,X(.>I!+E?0 
@E#2&D(BS.T;2RYL8$[.7(A)5U@N;;QKGY_ G.%S\6)  
@D6#S[4+253DQRQULG4B$[GV-00@VK-YF/([*6OIR']( 
@(T685K$A0:]")J/M="CWGZ.;)81)_VGO9P.0#[UY?.H 
@BG677URE1&X>X0WW6V[WN(V'YVE3T? 0R[5CD-WHU+H 
@"&,J<LI886="GFR35%:%FK@P4 F"E%AXV;S!Q9@MB1\ 
@,'XNW>?7A HY8;=>KS@65MKOS\O0]O8ZA08+*G!CP7, 
@3L:<RWJ+@N=BA<J7D>V"OY_V/E( NCDNS\L$4C5XWD\ 
@O3;.58.9^#(.O:\'>\^U" D*!L^_LT/AZ1M3Y6AQ! < 
@O;=0),9J58#P2A2(+*; 2VE-K$)@,ZW36 XND,''WK\ 
@DIH1#QJ9:(L"-+L76;4-IWF.B*U#PTC ]%'UEHQ1_EL 
@']WT>T2!;^Z9AF+]@K.QY4*;-9D+%I=/,*GUCXM[+5D 
@_REAHG;="_D\!X4 $IN:[;ENNSP"VHI:S[SC**0(LD$ 
@#'TFK]U*;B1,./'^\@U3C<0>"J?A)]&9>Q:.\B-1&M< 
@J[YA;YK+"*11M#0F)BAC"(YP:&?G*:9@'##(1K^8XL  
@&ABS_3$;YC$I3DZ346=JA)PTS7<TT+O$3DI.S\21<'8 
@]:G,7=12Q?><#Q/#$HI8K6*8%VLF3C(*RZA(C(=@C&\ 
@2*!_2)?8X/&H-ZT)_,MU6Q2_F\ILJDY6M"\<VZFEG*P 
@:=[LMGJD'' . S(I7^N>BSAN@<B&T'DYD.#6DI4G2-X 
@QA.=]F5#U6)>WZ$/8&S9H(O3'M%Z3N7%2!+XU6"WD9P 
@DHJ#W++.?->4A:):L=Q!*?F"YRRP6'Q0^8T:K5/>B?D 
@@/;"B9ZVU]4).,_@12H-^V[.N: JFK"N0E]$;C&];(T 
@[P!JKXTOA^V/676N<1OFF?O4%&TY3'H4/T8XA:>IJ@P 
@G^B3S2F>Z/Z/031T#^[+X5=TQ<".6XQ9-W>-U,H[>O8 
@M10P%9?P R& <\WO&*[->)J2U>"87" ;I+\;4OL7%-\ 
@$A.L5U"@!!+&U@4/LN<1D^.XV85W_54C%UD<3B(%HT\ 
@7M\F2*?'4WG&NSL^Q;G0F=V5P$['W53-E O3]1O2&)< 
@H67767#+;\VU,'M'N<;YR%Q5+"SJ,<\5_#"K4$7PV?H 
@D=M.E9D%GG,)1A?!IN2XE/'G9YB'L#/P]0]DH4NH?;H 
@$:MV\-^YFZ4KMMX+$=,R6:$\54HE/X$3VY )K8,DWX8 
@T_U;P2#P[1(?:=/1&[IG=OLOV?%L3FGMBH4385:  F8 
@J?--+:E"X$B.YB]F/!X*9ZBSDO!U4\<ZC4\P3(HT00X 
@<?CW@ZJL.]^E8F;/S:<]'*!;QH""F""X1:,CW^?=6=@ 
@H@0+?T1_Q!D4]D;FVPL(%1L!6^,(1JC3A]?F <Z<7+\ 
@0]#!G;(V5CX89-I?NVD:8ADK0\'KRGL;TT:'-DYMAH4 
@<$KJ$\ 8)HFY4T<CZUK*7Y]\;"N4YFP!F=H\CEWF<O@ 
@\F&M\T;2/.UCQ0>C#2_?.@;60V5; )8;?B\GBS4IC]\ 
@BV-2,GOP;P42CB0QKX/Y)N6+)W?$<ISBM=X;B1IPXYX 
@QA?@PVH+)A!+O6ZR*BTG=/)-Y=D7X)V2#CFW6IE9$T, 
@9>4Y2)$3YN:+ BVA= 3$6L;H*;#H1U2"0^C/&--.1.L 
@)LR4,GF>/<=SJ[?U3\G'*3.;I";_@TTC"G_1(][XWQ8 
@S*8@<4Q 7ZF'<&\U(2/A6OGZ8MY5PCTF33']C;"1RW4 
@S5Z+(TB3_D+!<IB6MM.&U#D#,;$P*U\*'G*4=3".$/( 
@<"<.(W[4!9OWXZRJ %B9)"-C?>GT ?BKTKLJ!#SG?LD 
@?>/!<9)2_<KZ8J5T<)&--6 00E>=^CVLI(<I1'J5O"X 
@CBBL&T\DOWSB&L>(DUHMTD4F9&S1P(IBFCI57MP'"SH 
@>RW><?(T>#60RZUET=KPV_5RT$80]>([]Z=\ ![J5FH 
@MDNN89%J1 (;Y% F%W 5XZ$BR@!<:E==\93$^:,3XQ8 
@D=M$P3=NMX]1Z4S?:6,"GZ5>V[7FNP6STA_'*2%8RNP 
@[&Y>*QRTA\E,UT.6ZC6G(SX]T%C%<'Z?&2L.-@*9Y0X 
@VQG64IA1]AHZG+#J1G1\EB,6)>_VLX(AB)I+[J0$TY$ 
@5]]&GJ#J[+)R;'*S &+<)?.41W@,\B_%YWWX@O(P)-L 
@#27^#\+# 2RNK^'T:IN8'1%>Z#TZ]2CKTRH3*QRR4VH 
@DU!$7P4SMZ<1A"0(2 L7;LJ+9001LT2+,I'3B36UZ'< 
0\\T(J5.NA965'*%P"</9!   
`pragma protect end_protected
