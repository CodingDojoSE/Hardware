// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 10:40:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DWTdNdG5TY1EVYVEDCuiIwUiMcdLm3oYsdN4YXvc5O9jYjf0rrw+3a5/Wsu+3htV
6FjqvwfJqn6C47Q9GebGgcI/nk7Q55LT2cqqY4wvFECn6nFgsrCtXl7EgqoPViRy
cu43YnU/dMnVu2xEApU/XQ8hx+JJxJV83JoW/YC4X2I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17120)
xoscWt5iswlIsn4Hw1SotMlYAv076ADvNEh2LsBFnZEI1/ZnM7Uiml7mXegg5Q8d
57tiHFB6qOxoaJjHmpJAQlkFTy1kPeO0qC+masXYnwFLR56oJGaMLYAkctcrYevU
0ggLWXzROa3GgkT/lLSHOCppfmfwtCx0lscPkIND3iqztm9B7SlEm9ROn1cGhK1r
qzK6Jx+IjkV0x9GM3o+ZVKL1LeMHraOEGsCujSEL4aNaFRZJSMBUmjdXHBGKZPo3
toB5l5waxsxi5GBSwXLExTahWkOdZ4257aBvUFYatJbyu6+9l8dap0onOXsY5rKO
V9Gj+Pa1Y/Ehv2XO7ZgMxPRh8GibCNbBksYCBBQYE3qQccmW+zaLdGlkICKjZ/Ut
T8nV/7Ge72fuKqkOQG6ay7RmfY3iNA9eSxVitABP6fm6ogPpEyMu0MX8iwzyI1QI
0z3SX/EJ97BNL1piXM7RKWaa48rshP05u1Ge/5x1AthKwS/w1kBrHK/6PDRouu+A
T+/k2mBmPulxep3w16AnaTpyCpMHQhCUxDWQk2RnZ2YVBy8ldQkSdDLc1QaYlztr
Has2A6iE86CVeGS4K9x0UdpESmtpWdwtVdciwu3tSuraGKvx0zl8As/S8JYrOFHt
9J7N6Y4/5MrtYpaweGN5Xm0Lq40bIxsrgmeKdnEoaW8fZoHbzUdjLWGPUX/cbg/z
DQwFfcpNTktconqumsRxAnVFTYb5mQalltcTXbU3kaZFOYjSN0b1pTOuReNBycBc
+SXcqZjMcJFU9K5WFWTUU0NtuCpVoU8k+zo+H564kaSHk5YWitgzbTOHcZjVF2gC
Gr1R9ma3SsQwd47g9m2AP5BRtqdlVRqnfIfw7GJmR37DV1yVsLIcjgliyNQGfSVq
iBhjn8cRLR9d57d4zPjci0A/eICxJgVrn/dDV0lKolRJyhCAHq+gb40wFG+eCcGY
FKQ8uQL8mHffeJiRE5/tnWaAl17DSQ+ah5pPjQLH2U/Y4ziVutlhbZwk/j14yt32
ln5acn+zrFQ4eRetuXjMo/6Y6va1pJIQcx9y9mVmfGht+2vnhR7P2hCbKpAfS0Pk
/ydzfHqYVlovlim3+gTKSdnHto5L0A3jmBZcel/WLAi+1bhwBIzI2PYndRXaSepO
tbAj6qsnEyB8RqsHqF6fNBGcBPSIa+wu3Dans+ibdw1e3Y2/AyJa/7uCvVncRAPf
h4UFRD65cTchV+6cQXzKigtwUoO0gVSaTZlsEIkBXs45oEeIhDehxv5SGWrxyQO+
7WXdIy24pt/fXH1fDqwEprKqWeQHCvRmUBCRRZ3Ua+YZJ7ssPngfq4y7FwcMnjuu
xrbPCiueqUjs8bdyBdVcU6/SgmRAFuVtP1da6AwmTqm/LFhMU8jHSXHXAGt+VDUn
v7g/+77ghqcvM2iTAiQD8rAg0cV5sIg7jwaLOdswymyEyNsTveEC/Y6or+/tHl4d
l525OyFK1P+botTevnbgg2/UdY/7ke62SNcG9yoSFYWZN9jAuvAby+KLCusCoto7
rHyNmivTobzSnG/0R4fIrS1NFnTOVjAhD1BY3oY3jvZvlXveCOOQu17GnzsQtD31
MguXayrjvNaX4CbnA+dRdfCc6S+M1xNYGc/Ug94xYZ9ThYVPD2iiYE8X/cLMGs0C
5l8nM+v09Fa4bDM3jMwo01lWqi2Zo1RFJN8anIMMlWBtC84BAbPO0KJTy0yLgVf+
C0osHHIMyN1Q9+ojHYZl9y26IKNqjVBmgFVNJqeG6+Mvo6yuPlRj+UgSPFoFzs1s
Ht5MGlB1D6QY7L4OK7K/t9+u9EtZdqrvFYz88eL5UkLgq7igJv+wjOAz7U37+kO4
u7Dlsx9eUG4dz+CdspAxjdjnhIYrtMKrec7cgvZjW0xYepLhxswL8j8gfu/OdqrA
q8L/TYRNz7V6podxNdQrjqWa/YxGMT6AxYqLAP6wPHdy89BWu98XM6yf9W3WK66v
CJnSM5IE6hU0Iw6RLkZ7/0Dp3TtHXSi1xq1VtiTRS5afaPi28v4eMhdeNzP4Zx3Z
2cjUbPIrzAo/7+3rFyAtgKVSxPKUhejIkmqIaZvL2E0OMLENMnvw2yo7Ta/0tkE2
oiahYf+9ZPT6ABwrXG4RXxj4GC0vppwTEIxkK3X+gWLU4OW2y3IksZB+oBH5+7lz
TqkSxJOZNrlDWVTm2deGqy0kGXLCWkkOcZXYNk7HsueboLW6Cw2Fr2MejGwFdCxs
8+JVOY8D5EFsMn4G1XwAdDAHIbKtvfVCqTNTB/qmAff80Ft80azOQo0kvmQbyMgV
+2LZAUOEmhcK4mZlMPqKNJHHsGXxIKbf9Q5CABk2Hbl7ZOavtNMbGBg4pJI5rKM+
ioib8kqx7cXuUfXIEiqJMvVg1kFug5drC3Ku6C/wtT8XrdEXxSdNqKpLh0GJ1A75
oLsEWbt+YA6/2xHoQjxH38Qw/bAH2wVWwibNDcg3gfvKUeflvpEd1rUd+F4UjqpV
6dGvmasZzfaVDXEzMpzeY1GWQd3CNaBQYBILrJbBBCJUjWm0o46LJ7+bbZ9nqWKK
OM6HMyYgzymptpIgcG7JQGftctcOO19cQaE+7LEaN6hhyjZSBcXXYjYDJ5dropPt
VF03hmVuBnnMHP76x+qD7bshbQ3rbGw3Zi+GVwtWcbblZoD8OqkW0mj8QGDsHCTO
35p1hm1vfGyqJWK6Cy8ESmFWGkbgE97PCGHN6AOZCEWcG0160AhgVSNtPxLSWqNF
WyJQEDyZDnYl+CTH7F++vzff0soFG03IO13CqzAmgbvDZ42Ie5H7UlzcUkMgPN+I
JxDyPksM+5KqWL8jNF4CPxleizq+M1QelE4ick9RiOlCYvo31pvx71X8X1mFZwvv
HhQg5u4/Ushy/Ec0kXLE9pjkXMpYoA2FqFxeL0b937QeyF187wPvzMlN8TJw2sXe
2Lq31MwYE8WJJsOKbLvKGMnYucP2AZ2FCAc4E7/OnezHq//afosTtOV8gNsXLgVd
gjs2nqmM46oOx1v4YqHjliO89kEhZB9BOg1TEi5lTKQijC2vv1Hf1kWi8n0t1dkF
fe/PcUshKyjTddEcFvZyXJmAV7KTdnOEHPyPaFVNKnjcdFSbI5c3rOjuurJycYLG
TIcu4Vsu3QEUSrxu1wWUo33CP6e6T57HkbE06bRhBgPnYBSeFl1bxTm8BNP3Gtyk
zAYDhJPFj4UunuRR2kgFupIqrd+3xT6EEhdesuR+GIJJIr/5cBeOpkOdfdUfDjap
MiTz7PzRelGT9a8GTlbSLYuGlHCKeDk3bu8UJBwhBdBP1ZJAYen7nG9koeM3HsYC
iNOdZUo4YIRvGXp5A2s6KcuzLlfV/a0uNy0xhAfkopSIVA3C58IdAC89nI96YGnd
6Dhr2Acq2o4Um8eC9C3lO6h0uhoJKzQx3x8DNaSii3xyotsX9ywzqZD6UpBzFUZC
EelcoJGsMo/ZaFfLop9yYZfWxdnjcjbnNfWsTMMYz69fZxiMD92FD7TPRHN9LypT
EHhdUCElcfxmkxaGYd+t0BhIQFd0DJYMm4GnZm77LmXpJPrEq+zu04CTmYiT/rRP
XixFPuo5TU++4BChhjETFvSTucvHlclguHpKXg6VD1id2XzRCthnOz5ry4tp14cF
fH6IZfruM6ORQdjf/4tAgXjKPbuM5Y3RQXpGZet5pBmft5k9TiX6XZiLREvheF31
pN5joB4YGjPyZyoGvH3o1IDDqeQ8ycFd6iLD6AEjZB5RKUiFSQyywuQAw6PYh0Wa
h6VL+My1OVz5eOZD/v5P3cIMf4cxCs3cPAI/4/oBNcgfjMT8BdSdEQBM0c2HY4Ol
0NpSyT13xlgBOJlfg8F+aCcdWalx01GFZBYv3qvhU3+HofQkE0DmiSrnZggKaP5/
eCSyo6jhBDKdXkgT0b8Z6q07NEjDri3W/GVb+9qNNZniXm4P/Nq753cOPVeZXsQ9
jrbhU2fhaYKrsDH5m2Sd5yNe8GwCUemiiN9YZYh0v8c1MJDek2aot6JC8159qvZy
bPCLvp2vQ6njV4SaZa+ootw5/gOH/4ZKdaLTW+8BgMWfSQdZHX6qhbg/PuN5aH/F
1XQ9SUCXyub73/TJzOywXAHoUwKrYQLGDBULBCx/xWZFekATjqKZRXZa5UelJMHj
CvlA7hSADHnB0NiT5xXd2S9fDVQrSoL+PH3zim5Hb2li4yzy5x73LmEy0u8lxrPT
isPfKflN3dzeLnqkrWEMpNMQrj5WD9GH0xslCPjAConvyVhY002GHt+8rSTCGIJP
VqeY1Vgm3E5oWSuSNYlHQ6KyneoPAbSMnNR3fIyT0Yi4UVngqKeXx+YjIc1vaEQw
zfchRz2aPap0DXiBOnHcFabepWEMziIDxKR0drc3+1w0TpZ6k9htfCcabo6YqYvf
aczVp98Sufh9ioo2YBYFIOu8DO8+9JK8tWGsgYY1RWmEOmGVtaPVWLFGcvI67EYi
ToBrij1LsKORmy3Tnfey9ox5WIbz3q8jEXCiiVZBjVwnvup1j9bxMol7M0kwUAyF
SkmDTcAWy/gK+9FsIpNzFe9Df6J4D80/lBOLq/t8+eZyUMfinDpw/Q5wFOWaFb3u
cwGZn4Pnl8ADKHYEtnfwVx9SqqSUk5rpPTS2TDgHrZg64+zzbhaFP2X8wOmLDQDr
x+/iuJvw5E3H7BHz+R4oOzyEOC6OPY7d0D3r+4ThONs+IZksLIfmkRDliHYzlO+A
xiJ3KnC/93JfkhJeOnbko9HewR5dZSLZBGsIPmKLyfrcPzUqo3HSuR5ygAuKgyOF
3slqsnr0zIrVtHxKYnsH6sr4go4gGkAJeWYf7zfqQZhpqBaqtbg9DcR5cb584jcg
GShzbAW7QIaK52bz/kdFKIhu046AdXsnaSp0yrNVY+CPzw0tZUot2n+TrtCOhSBo
wirOsHipjWJMJwp71o2bObFWtJcVUip0U3sPobnYoBQWiYo5Bs8021EWppFdwQLA
rhJ+fA1so70UgiBKikEpz57WlFw1xoTkqkCZauRmGXxzwKt/lPJCHe+4zU7MuZfE
hoPfmbn0ibCNzlaRXHDdtKbH5mB2HZF7p7rcgP0VS+OAoeCgnbBaLDxuJ1Jb6GIB
3ZjODyQ56Wbn7OBpOevu5bp2aEldXRc/9HFX6aQWteF41XKGfDyZGvIZ9SxAvdHf
WQXVC2odTTmaBwz5uYFOkGGHGl7gbnrsu/LW1YQ1hb6d9cYqoUTrsGZSegciD+E/
FFdsTcsY+dzSe8Cpb9bXWIxr18tUu5b7dma0+Do1qiRw3y/9GniswUQyMLw/2BOE
VoiFPf4EfRIUnkaJEN09CA9eFF2RtCHZxfo9whnSZ2n4KtchOhGVSHj4dH6D+FAx
8GpLlsVlDEvSW3di4nJETYB8oVJ/pYLmZlg666xh/qckneqvXj02S/5+Is3i2iZk
WWY6lGrWeUWyBSPA3phv5LUIMmtdQMLaFSdv3f4SjxN/OA9nxQ3wp3OgggCoMz3w
YjGZgBJuEMUxOHAoFZIt44zi4TCb3VQDRaeEYRNW8SeD8WCNnSTuOdF+bT9pBi1/
LsyCV5FikpwFHKT5Vi7rQ8VfP/IlMwGt5vavPz381DlWrwuA+oPA0pYbV2R5qrDJ
syjtX/dyEKHbTLynwHxZjLAo2/KHXsWU89Xk72Ytv9vcwmc7EzGb087BaTmLQAad
K+u0wpI9dLO8EFYinMjE0hwVj/lsdJn4SzULQM6p8evQuA5CWxuIYt2nlsp7/b+F
DPbZES5y78lwEncbxbhsrNK38Zhb7uNjnKFVdiUCIHBy7xd8yt/epVEEND48GGbd
NqyGCV5wF/pIjPNg3RtaXqCDEnSR5ft14AkZlyvQl+Ndjz7Zx8vvptbvkplpMgt3
UcC+VaJ2IPpnueHKzyxeIKrlTzWWVMZLX2/NTa6p11MN7eZ0PLdkZTXjyQuhn3PD
JN8YaYAm0QfVJcvypzhW+6BsMNBJVPt6nqyJwEWVjq2cG/XlHNN3P6csv2o9UCpt
IruUvsH3/BiCHu2QqnK7xZW6uw/0LQnX2qE4a4Uysk/OYgt09Q8sZ5YnyZS2H7zF
Wa0nL6WjsxGeUmdyZoncXfPq9EYsCTRdfa03An352ToHnQ65WhdDMgJfrnhL6UFE
6QjR+2Y9v/AUX94YcUtKmSdhf8ozibvC/NGicB4hHnueKTchVg5eFPlyB/iApm9n
1FTXwzYiZAVEv4d2S6Or1As8iE0Y0UYPnhFX1E7fgtcJw38Pb6xEdLmV25FXuJeX
9dSCasIZCfkdZs9pEJ42G2IJJNPk4YV3tAwLpJ/l7kHgMbfDTqMACYyJ52entI4r
qZa+tT8K5da7ZMt7WddDlwayKKK1wt/9UR6Oo3IWxALHt7RyGJ/f+yF17UB7oEr9
hfy8oWIzjzn3O9UdmRGKufz2Zp0pMh2zoeC0SReplSSpSnweFC5jAM1mqkxh1NXt
egiI5Ve0wnBaHflWiiZBxJ8lM1tCtBwD25iZM6kxo7CoITgb7K2DPFrONbSI/ehr
gcqGIho8S8j5GaJnhMj7M8heDqchK2hCuGvid480sKwC3dYMzB7vSlM0NoPH9/cW
juI0ygJAMqjIcZOQ0j/Znbi2kwgiJ5h5tE1mdIxWZgO8x+0Jn069qp0BA2ggeUhO
G7STcoC+95Gc6DX71vdWOr805PN3uueQmQYtHGySPdKXLUYR+jUiJbuftxlszl82
M0/F6jwXkudzXSdB2n3fV0qIyuo6KgRsN1PUtr8SrPRUkQD8Czeed3iUeKj1ctyE
uDnH6Fdfn02lUh77GkkfZG8r8We0huITppmSQ/QqHdifuMgKqjLxIE5eI1twaQ/R
0LK7haj/JVXqhiZmv0h/bQtuaaRHXYapdmsfRE1e6Fxy+vYZXe6shTR8c9tE8T52
sS/9GLxJRH1zqbBjA88V/p2j9iIcO++P0N8UZgUXMmyFPLfQjPfEWDFq8MRcGkwv
1DNwxHOKXn8FY9V3njQ4rEiOXDxI/ueI3Akk/2EkK9PTA1uJackFOdjUDm+fp1CG
lNeCRg+Sr/FXfYHn0GHt1YaWyT8smC+W68RMdjhvWE1UI2HIsaMawmCEcBl+e1qM
p4WYlQlkvbQfc/WjSK/+SJ+D5EKoyjVO6Uh3+WYne79KNRfAIAFVkx1mtvpas6AQ
USMH9+mfmdx/mmCg+TCQoN7tUeM+JBx+lM5oUJ2pM5umV1mQD2UyrzfirJrPHknF
PUW96XPzDdc94nKbm63EdNSrpLckXv+CsCHCWWKZ5w55xJOVBEdzsI+m3duP7rvA
oVUgtRJFLn4XOM1eCtcrXcYv8lAAMRuiMZcrnVlzJEAS79Ug9I1sJx0urQbD6a12
jsp6K88BHdgoEx8pCow6VUrsuU9OBTW6SuqT0WSZjex8hrZecDCeS60Carbb4UAt
mMS+W4ukytrAEj7Kk0np/9BPZPbMps1lg/n3vXXq0LN7X0GxyjVKDrtLIOPlTDPV
aVIR6c/OMfTsYnwubtT8WyUqOZyWSYj2RHeJYuQ8W1TM9iCjaQrLfMapWcFBS92O
cJeIbhGbgpktGAB4F/OrzeUQ+S9H1YGBQfunzUM0l3qrlsaxRrpMS94/p69mGLHv
NXjvQD+VrjLb4JSeNgjisdeL/+GPXLnJsdbInC0MrQVGdLnSVLk+YJmpcx5be56U
ai4eH0Y9v5S9I/YM50BDLDn3T4CQWHLZbCDRpBXoksmSJPPA8zFFRtZc5S0G8JKM
HqaivoN1rosTZccK+gv8lkrCcK6fcHkUp60/sNIaQDnkFBR++4rK9a6O1T9IWDO/
lKAOO81WiIK49HqyLUf5uDRPGQlS0VDIo4WdCXDXym6u7COWzWJdle49N2zynPx1
nVtqd9ax7qeq49W641alUVYFlDrh7/GG3AtCrnxwmXq1gNq6mg52hHPpB78l6pQy
U3hryQPHaAsdJhk9W33PDxh9Tl3lDVi25FAy9evoa013U+2j8IOchiN92JkW1fYX
Fvxp9LAWgHRa7O02+dgilRWVUU9lFBCgmc5YGvlMf41lpVUfParf3twzUR95LR5h
ArH3PopemMW6IPFpqnYll3w2hjj0Yt4X5/AcSZV7dHUbf26G4XyhrLl8Nb5P9LAX
/4BY/nO4TT6+DZZtirMr/gBNByTReqnkJjRDkMqLHu5kVB1FLrMbS/4ktR215dtb
xyM1MYtcjr5yoI9i66ohSv+9v1haR7l10pNMK7dF+GDQmKrvcfWm7R9liHCnMg0u
wiI5MQeR2kZL5TRw7W3luAwrMU8Ha4QM1Wml41a7VYT9IPLv8QtXjcCz78fyNBOK
LFdBVsYf7ujVG+xSxchREO+HYD3kev0s3/rQubCJdGpmkYLSSTt1klkCgcRLxhLb
CaoX3KTWrhCY+0PxdgyiH5Ogic4XMwdMzgjeQVTnV9jLcD6Jz9cs7cXZic+aIsgE
yaN5usJQx+BXOdiuTx2zYpbXmgxpqDXR7X3rd0nGFFUw5wwYHfhu+6EUWGDKZqFj
fsQBEnO7eS03uAu/Xh39GTGybUBwGeKQ4eNpd4uepUreAMBpfCDMFmRwC72x1PFa
B8zs/oIZnmPhHhRAfzdvSwwKK38unfMTLhZZ0mBs39mBGSRMsx+5oVwYzY5Sv242
0OersHns6cOzF75bntvmH027WE9aHsc8qVkcUDxY3jd665Dngx/Q6V4yvdh92JUz
Xtj5GgI+HTyXIoQUcJeLrkHq2Z0RYYyRH/j/no5npxrASBD2Tb/6VUws3in4GzgI
Fs3LTbalFqlzamte2THLxWz1aPGrkByESbmdi7Sgw/83jfWCkII9GUm3O4/4c8AA
0ZKdfbnyaaemMqIfnXl5dbHH1+4nZsH3yoP0Yqka/BhBTwz1KgZ/YxT0lH1Isgzs
7xNpnrYrYnl/1kL56/stkL2ryfIRSJDMg9LIGXPdUVPNJu7pHszmpyfozKqhwgMp
ydksV+GFCSLlLYO4c91WDGv2Rjvp6S8i8jmXGClyW/sNJZ0TZ8HgRu2AS4g7bBL1
yUQWb35tPbhaWGh1TlP9hM6tcMvUNq2DCVp4IVJygdKHv19GWrX1kxTJIcofOtAp
bGW2rHlJJ++BnHC/UuHjkMVU8RTYIreEIsewHOWw8peEPBYEWFoEdAGHjt5L7cS7
5QNJTnsSwXLUufnuA/fNefRVTF5OOUoI57g72X4+SQ33XAK4LmoBe265zpjP84Go
AVFdj5kfzha9sAvMCl5SDnGEUAcgwf53T+xwhIzoCcIFp2wFPDue+xUjRpUC8cjy
ko0ss41E/2Ii6k/BmmpHWyNAnO+xRRkqljrmIkyF1ch/P2v8EysKdQVslOKfZHZZ
ckc9fsbVsruErkOCDjdOKQfTqob4MJY2X6Cb7coTMmv44Bxkw8D9gOKOj59E27EZ
SzJ2eq1O5VsPGXZ6rf39qKEiLpU25+TAtokxNOCfNgIcjBErTgUm7TUusbXZnM7Q
9ZiSaURkmXimCvDxnNCjSP/fCxIFXVCO4i5cS3pVMOYOrMH2+c5f3P61C0TMfB+f
aKXfLIVeRNRNS8pxaWZrvNb8MxOekhUzRP7XwNqZwQmxLFM3BRFbz5PKGcv+7avw
ce7niP+sX4NSmNfBmND4phpB1KW9vE6IIRuQ2md8LHb8rXE5dB2kT0MnJ0cIfBYN
4BEz9na9E+ojOjApZZrpjlVuhCQKeZBTk65FA3WhtJLGuf6tf6nwlACsRHxUrox6
qbbc4p4A850SCYdgHSlIV0qAJnCZQ85feBLzdGh8G1a0NgMhKSv1qzQQriauOHu8
/NYbp5oRELa6jcM5vY+vRhtsPqnOr8CEj21KTa68PjQt3jfObVjLiJOmhlpjAMmg
/zQE2/nSHQ1MwFgn885JS9ACJjUUX7dooaYmFAPwU+r45Ms8V5Wnex6gIDjjqQFQ
xW52SaNnfDNoKf3WKQ8802oTN2WfkqSZGt1JGLqF4hO0Ss1WIDQoef37ZYtgDPzL
ERXhrVRJs2r6J1xndIMUEn68gCniIeS+ZSQoBJBJPcpG/7ZElwuJG8R874ujJrXZ
KiR+xxlWkEuiSJQFJHqTbNhEJpE712ZDihzoxaqvXGuCFhsJ+oPcFkn6EBzXu9sg
acPrLL2po+AKgygxLMEyCBSKbqlUPLCt4zNT+Dbt170yAF7ezSn8S89o5ith8vzC
57QZR3/YNWfFjU6zISBemtkloWKBn3x1uGm3ajnowdtO3fDEWOiXWlZCI6M+7U2M
3ZchCYuoLUfjKbRyd5aaIkQhcyTa9I8kt9765GaqFmi/2+eW9Q7vA1/FY5pXHHnX
zW4oGaGUW022WlFfSAQZJazpLjJBPHf6RZENgGTgHGTBepnucMDBYEvaYV3eUbWW
wC38Gaw1LqXSG8cYW2H5vzySFG7NzMkPHLQ/9lwPzwUZescHPyDKrdLO3BJsZe4U
SXAIqMnsrNaSnuB8pRaWV2xrgs+7vAO/aVDsUUxt+oGYkvqXBUE07KEYc0g156CI
C7Z15RUHoW5caVLqwN/ZOPWqvjLEl4vGcSFzBTZl1HOW1dUeqwctzRAJFZ3pJn1l
IqyJNQKBR2WZMEeUv+vi6YLwb+ChcayXpXlr9GMKfET7QCmXL/tYw32SpOCZ6tBa
nXgTFGmzrugg4WfjAedNIFRr8AUlW3DElorEanHsUX4tYhlSWwc42nEwCobc+lmS
3FSg2hM0sLO3/aDVjuRv1mUy79Nj+dYsSY8i7/9cxdMl5C6RJBvVDcpVxudayhiF
zrOxMdXZEh74AvWWuS8tOuOJ2DIASG6rFioKSSrEajvvdWoh4kAy63VdBzDnGQWA
sFkf6OMbmSYcJ/ozBFRyxXqzn3+upFKhkSOI9zWf25A2mVVRDBmYuM2jj1fhRsEM
r5DNzejQlpjE73q2dv7Dd7ex24IgvV9kq9J1dRPvSou5mEoTZcVHzwZsf7Zs4hqA
BxlfTXCvDLQSVAIxajw0VL9oKeFL0GG9QKkt17y3qdIzHCeD8rpiFECowBLUE330
AZf609p0V8CNxqfwvtNIOfD4j/nYx46fRlpu6Ge/3oqT2FwXBYWCqZz7doosWqY/
CeGck0jKXm453uo+YoMsswz3og/giBiIJuWk6Z+Nue+2rLwcpmDX7b2Hcdfa5qu0
Cre4MN5MEdFhelTi1LOmMNASg/eo7fpndfygNmFzPNy0iCZPDfD92dYdrFx4afag
uM1N4OvpbyqeuBYLX4R55X1NgOehn80WL7cVTbEcge1hVB6sHLx8khcQCzJoa9xz
gv/0Uo87zYMLOYXVaHBobTmKsfPYO5srEVNmf/0TWjOQfrfq3ZI9WQRMdVXXmqUV
1DOQThZkFBukipB3ZmIDlgUzcX0W2B5H0Kn8E2H7bSor6lXUZeRS92fIqww6wSMm
YGDQzgXDSwFO+HzOHytMhtnhF8p0rLzyw+wAOoGYv7T65wS7HRQq6pQ8iYxX/dD1
pXPY9jSQ4z3frLQ+klL4tcb5OAQ1eeQhSnZj/+aqWfG4bMjAmRDlESq364dtolML
pD8WCtWRx2WUFQq4U+I1PQStnr+iXREIoBxhwujZPobJv0KdJPHI9txac09Aw/OC
w3NRZ7F9sAEMi0s5PLzjZ0xw4K0ae9ZNIzFTWeVSIMa/ENm+0ScsmR6LOYT58qOg
jPpCn0T8ox8jKQ9Z23Ca7TmpyO8dQllf3SsAgYsuDnWKcORgCW70I7hdd8iv4/I3
cWJ+HBPEIFz2uNF5/NfmJODBSkTnuOQAQYPA37QkYIyXv3LQL2Y6icx9TUTtlQUV
06ALwlZzu3soz1NYH7I0oTGZNmtNOZYRv7yhSwavRr/6GQiWOYZdmjbkW+FgHgiE
mfvm1UFpge2M63ekqpUAu4DH0xFFggdWwzat9YjNUaz10etvyYhw4L0BehNVZbe8
QYYSrvJpCUp1yidlKR7iLk6XoajaTWLm6E1+XTOhdnyeX5jTQjJ4ygl1APo2jnRW
Iz10ZLhap4T1P4MxboD+qAAGjjBbuMgX4OZFZ7v9zcYtEXfyEQAz7V1G57e38wL3
AJx6hkDepuATZYmicoNOQD6G+TkymLOriIoxNCldVN0V6clujcBV2CUm8TvzxPR/
F66tRgtkSprjwlqrOVoBixizE7VYcPpoNMp82O5IJbt7e9g/HIjcpHsrWlQko9a2
VuLgaE41j9HGm3+ZxhzR7xxQt4lewEOWvjj1RH6qMPnEgrI/DvVOqqadCCGy/h0l
+geqNo2Jhgf7s4BZizxg4F0/TwuwyysllMrujpgpovFBgmB+IVOnO/NMN+z/iB7I
mJQs0Ux685ovVx9Gb8g1IItiAhIhVavMqwQqBxMsDNJ4Qt5pnv4C9WoifoaufhMp
OFopcLLd5iwjhXTVU6POOQB2ytqQMbOIrEcB2lF8RJvbrBQViuDUmLBoRqpmG8bD
BMYl6mr2NqcBg4o4Pl9XxyXtwRu5zxLBCQzjMCzrrBC2iohniQHtSRwGYKwsU9Gj
f93eKkJuH1O2ho6jCgeSWx9CTDJHENrf9ugn+fTfopPDnZrV0QdZg+hoV0HgMGug
d6nR1zoscrUuDRggcZ53My/Wqepf38Dgvldmi6dfRWz2PAoVs5EEg/6ELRH8F1Y7
BAs3dBGdaAcrZXyiZsfUaRQmp0pYVqTIV/LENLLtDPLwMga2LoMpoJUvhhxY76cZ
fbxC4880OCNof8Jnlq6h3tSFTRoflCV1CIQ2lRdbnRXtWZWe0UpEt7jG0iJnZGN/
Rh7MG8UQZzqRmEnC/leTrcduI/oHMhtpWkZ4t/wW28UqtuFUelTlziLaBr94amqO
D8IKuZUVhV+PGi/MwaEBu9L6D/dof0fwDaEowXSEcBXrb3y2rOSu68mwAVDjEKtC
M0QjAGGJaht1lRWzDlum4mpDP9kioczOh3o03n2KTpBakGjMYYQyHMd/Ovltqhyi
fEEmeWy5C7k7JeE/oWc8MOiWTeG581Yvy7UGMbOHRY949AXJxcHNOer0zSNJVVW6
ZxWOLQqHcwDixHD0R2/HJjexk4HPT2OjZ7gUm+yU9qStTErN0863U51cAyiJlCNa
hYy6sfL8QByRVyL/eXEM1+KrQeTX4yaszBDcGahViTk5upigx5K6GvdRy7uhIrlu
EDuNKX5zGxMoNKzHnQTlI/VPNzwLPByj9jDsrDi7MONhbEc0P9M2YZ4oUX6t05hf
Xk/4yMFSTXXqDNm2mCMsZMYz4UI5TVyDoA7S+zY6yRnppKY2ffbtfD1tx1ptKvyZ
ngIrVLirjj180owz1+s9xqFQyO0XFtNtJNCn6v7qRh+b5LnQ6225U7U23oL/wtxC
FHCeleKLqlg3mCqUPPDZT+hZY26K8ZCXDXwc/R4ghs3uinRrESiWdVxUSDXabOuB
ymx94VhHe/IKi2IGBsXvcsIQffuXdg7Lb1nPspIGJqm5xaszWxCkn5cKej8khJyz
jjUWQmaN7P560+1JqDXDUaAEQeKZ0T0of4sm6Niyd98MRguVZOKYUf2923fkyJYM
Vz0E2ADdKzP99+AI9yYOMRc37wEEV85bEey8S7IJRwGMW8YwLODWHVsAmy4Chd7y
fQknXK9kGXqxrcGobY3Z8XdWIdRZPzTjMZ2haS3x0Zl40Td5bythDlu+0zklLJos
oCCjvNu5AzoVo+h2/3WtXxTi6Gr/fXVu86MExTAXsUYTmIp7MITlYQmgsgPOdTYb
oGtzCky/+LvuDuJs2Wur7ROaIRjF3P3KB1T10gUYHSX13zcF4HFLyEVDjPP3OD1m
4ZX9WgGEhmxRn3Ux0SHplCff9HxRAejn58C5whAnNAO2I8SRWhYfuhDzz9apkDw1
QoRD6Vk76q4tYQltSlatZfbssaNb9aNmZoAJNZRLbLmZ2zBLmBrM27CBF3E65PFH
Ih0wLGM5Zz6ByVHl7y4/AQZvVFpHTm7/mJ2sNd3QaISkDqyfZGXW2SBlJqEd/Dn3
k4k8icrlf34TIDrj9hbc2fV0tueZQRENfN9dMZ5CJ7n3N7jfDib6B1hqfm0zZj6/
QCjIqDF4PkiTUpb2vTuCLjTGh+ehmdwvPhaIjdWqErsb0pdGh4A09CnrZUMOytoJ
aN4qgQ9OD/acconqU2hmAsBoGyAXkn62A6L6MZUfGKA1ixh9M9+i99q9fsVpCm4L
IJnhqF+r1NwCO022SDsuGGcQfOT/NsT0fM5iQo7Cs+BPujIerXGvW/hhGhOQ0y3Z
1Shg9Wx1hqFVHfYJSIuGLzxPOrSJVZfoVhExW795xMbpXQz8tL4AE57H2LPvBahg
Pqq0DLjV3vj+0RXVf1WFv0a9NPFeuxKCnlTdkyVTiiIQZ4Zw5O1RBYJV3n8hU0FK
i5oj3XiB3LChl97rHCsJ1EwVkKECr1CK10RgfAQvHwdfDwZZ/laQwmzZNuMIBvbN
ZUVCvRamWVcBEjSOJhKwbsV1L4Bx+jMRzqYvN9aCU1E7ON00h6DpKiaXuQ0+6sJ6
JqJ/MPr4AU3TsiRT7Hdh3E2c5z8nGWjSOzIoSh5LAF8wCnYQFfK6GDJwmQp9PiaN
yWSEiFzSD6yN0o1gRg4zW/B5uQq8fqZtVvsZhM6MrmwnFASrVz49YD6AvDD7HfFL
J7PSUo15Xjh6ya53Ay/mgVcKktrNOh+QLmfZT8NshtWUwow8+AiGpyOzIt68Urk+
Uyl9r3jl9cLjaSrlOA6pVOVuw0Wj4vwDghU0vABXJOtkzWUoHFeLN4U6i0oOK24L
MSxv0Q1RbAoS6PQmShojjCPo4Et5wTIjsyZn6WxNF98GaShxAaQ3NizpkDLbcqtg
BmMABL+pMK5fkozSIzGorR0VkXLBfCpRoGQhO2JpAO3xMNxtg9l02AKWuga4iu2l
quZqBFK4YcKbsToMXhlyP9EWIvQPMSE9iihYmDQ9zgZrN8wqNgD/dsB1lT4aSJAu
ChrNnd5QuDzz4UGFcGpKlp2F/EGifUfdy+JMTP500iP4sMlHVQPi4DmtDEORkVAB
aQbzyygJeDqDppBkltJhU+0k/v4yV60Pg9+vot39omEbEX0EeXjW6in5aup4tGSE
dbd8pFl6K0AKHgCDzE047VPpKD0D2H1O3wvH5SAZKGU1y3o+dxQDRkoO3BuWfryx
6hrS0NiSkeSBhjQIhSscnjt66CbryQNYs1VMlCSMFWlAaVgOtZTNv1Y4COuxPfdh
wJrwo51O3Il6tpYH2mTAKSRnenfLMsJtAMGO++eII+Tz7Viy4mVa7OIf4G0d1Xpa
w7LVqMKH1w7/I1Cs8mgdFRePYhKMHSqmzrXHvqh8iYLgrGamAmhlfZd8fOg/qPGz
sS/VjZroiW7KYfx5FPC9LSl7fPiheNeIBth/RlqMdvyv+qA9rBLe2fyJVbG74jNy
0DWqPo78FQZDSRImvNqFvXDCdZSpDlFCgXo8rP3RoovOUWBqIU/3vSUO8w2KAd3S
vzdHzqWWHtyrGL2ciQ57fqe6ZMg/4Q6m8h6DMe8iqK+Crk6pRM7HSLZtAc8q2vTG
Awvu0yS6SkUpLZedWrAEpFvwfP5B3mHDB0xwlp85erWCWyY3eYv55Dz7sRy3DPz7
ATniYSoLOJC/mCrsEmkVIp0dzvdo32vgcwS9gRPsKw5p58DVxkCTeNiNYoo1bTWA
M9WhREhGL/hsVFRx77YptURZBL3oOM5BE/IuDeAXMGj6zOZmTC2FsU6duZEvhIHf
IQuPgelXZZk295uFk/HcoVP5NlbQJB00ny3Dux7RmwdRFIkf85cfBhBdSRg4xUnt
zwL+blJ+Gr52JAzrgRb/radS06Ohxye2kv3n3YOB3HZ7gO1jQ59PwrH6rqn82LOn
nAkAMKyMa8UUPWe7otnmz62xTkUEmH0NBsJYTBPqD3LNWrwezqAHzlUUJDukMXte
cw4hg6UPvugRfFT/9XNODuy7MwvdGFBDsFwfS+d+kUIr5jTusuoiGHwUERg1Rz3D
OxvQ5/PYc+hdzrXpUHzTkm3LWBpxpLfoSCg7tq06roX+OjQ7AX0TgovTtj6iIYC5
aVqgWeBgD6sqmo01GDFgoC4QG3xyCgUdXbfx4fs3M94kGRXe5JK6WEPS3/Vxo0Mn
OpCNMZRisBceqVEIkEEwuoAVv/aXqDamEBww1tM5h9Zr2qG4VfEJzfH0C68ja7W+
TLyXEqhXV/MTuBGk/LjRUR6xHS4E4PxJIIARdh6XuurUmM5DwJ1xBtD+MInO8LGa
N52hFyI3pG3+YgqB4owP3R4FC9680JyMft4V1a1PvZ3niqFTmB9E9Br+dL3nBP49
qNIFkHO7iml13Duj/RDO2JelPF0g3szAkfQqCsdXbpnsKX3J6kH+ynq+nqFssqZ0
iVxXDEAFlv9lDe3Uhm5qEIyCWuN5F2zJcJIf6KPbkV8zo5uhCVpfomxVCajbGnGR
EnDIGNqEQEd9FUWsWUYl6e59B8R7p5InWTcZpUJDxLU9cRHC9LCDoH2cJ+/3k3oz
j4WsoeDE+dbxPg6m8tJvm37a5WbIgAF/KIY572+louPIff7TsxmrnvNb8TnBhI5l
/cU8lviLVG2Vx6HrMUjXqRDg3/tTGrglKbLjlGUXE3ThmHrFYovvX4SABtK3fmZj
jpx4wvxzC7aKI63K751aXX9xvslunB53qHEDdzsG6z5LiE9tetWjnAU2qadqboNA
K2Vd3bBSz8eWJQEtNcgiN+THi3PFQ1sZh0lT0unpSlDkvc+QMzah6baqom0hmO4h
m1rflqkxd98K6rKjPIBEUgIwKpLbfu8ubONKfKBkKnmZxiG75BljPRSghN7sw1G0
fWCKRKuTySJf62YI3mFRUaNQ9hO42GmHg0klWoiadH2ZZtrTejmgoLw4iYNEPXQc
qzb5l56DxoljbBD4zk35Y0tTvckghSt9eGtju8y328y9XiC0bomfoxSxN6chhT3M
Q3FYLqEHWRpjPcXdUhI72LTLJ7uynavJin5kHTcrofq6lAoatbv7RU2zBuMt+ALQ
nuV1Y6NSvLbWCUKUyFALeEENGZQ3s83JtDc3nicBeugjqqenrJqxH7JIDbgi0M+T
T1nXclFonwoYJ5yB0qsT/ESp1bsmBe4AEQQJFuilQU33yKNVSGlOBSAs09uGDX3/
VNcMJR0YvamikBRlIjUb2ohUTQOo1NvYaKqyXfNY2Sezy34oFoVx6T04u0qXVc7M
MO5NUMfE2pWvcpdXI/Ef1r/hndDmqH/d6cCjDkQxUj6veZ5BEDflHSD0YwLdVbvB
u8Xkp2Fma58WFgMdnxaszAFGibQ7I3Ylhw1l4ZqHCv43t4HVwgcVxXl7YLkCpYle
VlFAdViRTVDW77lwBGCauBM8GF5bFbLNBaN/9aWkIx0JABofA4ZVuWkHC2iKkL7P
ezqvvEFVwF1zqY+qs9WAF6qAY+ofyMemzm+Ur2Rz1csZzT7BUflmwLIYPf4i9nqO
reS4WrZsP5wHbu2Qz02KRBlayjqk5LvsFdRtMFh6srJhzi96QFomn4VqIdUocz/A
Rjv65vAYLFL3CMVytvqH2gFdYml+4VQBiQsbWC5/L1XrJXH9E7bG11xv4tMYhiZo
yA/LpYN8++uob9qxUZH7hX5f4JC0Ol72H6vHzY+awbgTHmZ9EVtYAdSwGlP0q18C
YtQNkLgWPMhFQLXTHL96eklUuPPxxD7lKUqOcYAzgmGXWHqHPy7Cq06Vz4yJjiKe
OonGvP+ydYfJDiAed5Ye5OanY2jkSnqveL002WdDcESUxY2xmLQZIQy9YH5LGpX1
spAfL7H2mGmWGVFkf0071w3xxcumxTR3Mo8rDTN/+eulAMFml1KwkaEbJIVdKVMZ
9QklfWwExRsjGj1mL4i76Sy7+ALgRN3G98lRb6HaqU1aPFc53v/BWiUA896nXNKu
oH3YuLv0gY1NswnfTeIn/BVD+dzMCqhpeOmJ5LQilq9MsZaF6R82ZIVcFnyRUPK1
t4VVQM7ImVmJ09/uP6QfXZvpzDAm2mIVcKm/jPhkD/ghYEZFzHb67jkpqawHpWfJ
dZMqcbCSDLtNGAYDvHF/4HhWGLZWSy86D6Iu6OxI9kXLZWTJ/m2DcxB22MXveu/5
stKvy8LvQ2gTWneSQ+mwPK6CObUsT3/5RoqHdqyAoTnDLSE000PsyrXkTijoyHaV
Jbo3TL2W6ZV+R7EaCOeFHiEgrD/4r5D+MmO9eYZ0m7GZ9X0Rg5VAz63V6ZEJ+8e/
Y6x8uFKANLT4bKWL+jirWXM2ADuG1y7XcCOdtF7jhaYEqGckT/7I+uWNXdQSVk7j
33fJKa3lCpkfQLQIicEmKbhmnJeTQvvS+6phkLdRvBpx4MrG++ZAUsosaPOI3rvq
QSZ+zpRColPgWa6Qnq3pwVUYSYZQqEknlJrzomuSunBqm9X2yUo9MnxezxhFoKJy
KqP56Z4xGK1ICpFCBtHEZZugK8JbYx2o0gxiVqtB1776ZpLLKic9mFH6LjPToQUU
+Aq7d4bKeNWWx6qJN5ZCrwcogcol2WJ6ZVdB1mJuq6n/MjWhPKxLgJkPnUXL9OIK
5idna2E4M2k/PO7Zntsqc8Rpkn9xJMVfoSyV5foxtJH80vDzA/hOv5Ho4a186yqB
fUfxReth+mlYiOvlcOFRAl/Jv8PjzJ8k7A2VkLFMMTwLA8ma4GROXurYaL333aso
5yAPp+4dQZOUiIWx/CJbKhWGdU8GcwwA+KM5pL27dubzYaLssPiQMBG0zGtjlvMm
Z3+vl44qIMiFEY4LKgOfZuXy0Jp4VkZ3sMCgQY6I0x5ScMVxlEFFuyUBwgS0W+8U
YGOxBfOccibuyCJMm84015X2znz3eRnJkgMQ2saxOZAc1d79mKRAYwgqV3EsVPTw
c+RPX+mcUnePiQIh048hW24RtU9cZXB6NLWLS+1lSXKmWfNbxLRz6jp1hg2G3eXO
Jlp2eg4wL/d0ylO8tKBZVgyJ96dpd0PFQCrRg0i81lMq8G+8RfKVfom+HKDMqe4u
1gom2HrU8MhBfJczgCa6nw0jvTv305RPVSwLgIrqO5OFkMBmg5j7O8rhXp6b9G1P
QPfAulKV3E7oTRMhrqz5Xb8W8n7n0mXXjPFCdpk76HgHyCt4hay695W5ZaMCSf+Z
/arAXvAppu+3BJLw9LPeAiPYyhuAeqJu+iQSe1xrQ8iyKdkbDAbgylJQ/7+Io+MT
/aAmWC47ykVJgqHsvflMTbbx6pwv0ARukGhgvoRhlhSOCRzxHr/xWz2q+4XPc2k4
fpCEpzRsMw4/h5sopZNAuoW+WyHn6fzToD6ePBqqn55xsJD9a6spf6CnSp8Hj+p+
z2/aUIb1q9boGlcmxvZbbSy+LJUiZJ2McDX4sjvqFQ/a3eq3mGDpAgTdKB+Cp4rU
AP81c4Mzp7kvng2tbDs+0ZUPjByhQ+YXAnmGY4vz07CwVv9ueTvh5ML/2Q2VNNhn
sCMLf/bf6bLNv+cbn8VJGslB/M/iScni+TfeC85YZGDbC0zHQoZAfQlOu8WyPPu5
+mESHj+/6xxu1WQkjwb4A0WiPK7YqlT5rH26A+W5T04+4MYtKbDMZ/GV2VLNEqCn
EluimebXVqznI9kUf6v/GOy07GcjnmPclVyfjANhImuOcsVVvZl6c6W6nEAX9c0W
wXwgsIGcDXSHVe/mUwNGJohaE3LzjQat8wVJVcto9vLYGcb+cOYIjJO8xWjvkNk4
r2lNGMF+pkr/RzziPBW/W0CJlHI9ZDfJWPorQXK8ls0p9OSFhty7bOaKdVoVmd6L
eE+UvNLF+oM2wtqil4xWiQURd9dkj6XQM0Xcw7ZMgrSxMyhb42yXJYhO02eVjVHT
Iti8hHJBSWNpm5qEucoYsyzDMlIMlNxyPSFgEZhA+gRUfG7jY+W7GSjP9lIr8H5/
oMaEkK2U7j3UyGYZyMMcJ4w+BWvwVJiOogpEchhx4Vh++2xvS7DX/LDKwuyki4A2
GdJXF7uEd+lPP7i24q+EoZPIxWw0tZGOLwfCOcY6MklEkVSqdirOH2eXbxHFIC4P
k4LWja0ZsDm3prT4ZBvuU5oAF22mFJ6wSEEnxqvuqUe3haSw1MuAv82Yxhwjf7ae
nchkPTrW1QmOqQOzcE6VgDozDtzd8ie2isiElD6GjdR1ntGXbIpMI/GspE6GcFKu
gtRKI2aKH20HwJCljIjQ1CM99KQJMDdPuB2KU/x2fAmJwerl0f/T3IDXbfgmr8rS
7okcrl4nufGkoBs/TqBhxdEcgmaTtYR+nU1lUK6VzedPQfQv6jbkMWACvQGuWHtv
B1mQKRxH9O4EykKCLv7tDC/F9qlyv165kjUzhv0HIdoTRlmBfbsCN9ZBz3KSFH1k
bUro4gCETN+6+pEqMjwCJpB2qw8xSVJuH909cbzxR/AFNzxsBKDexiuXz8FRQ1B7
d8HLnTXE4OlptilJ8CWk4q8tDZscgbBgGX0UcdfQ5GGsrnFuy5zeqqQbhfTc597L
Ae9XwfgdeEGl2CA+uVFh+s/3d2POwjuXEuGgCq7VysA9MtKaz/3Pl2fHnhq4Vmts
rleH99xuPqMeZ97ETNK5585h71SM43FOJivpcQiLHK6xWnxZMXw9bxU6i6thqdWS
B/tGISb9594sCYnRC4aqpYjmgRtZ/u66HgGuz2PP0aeyqZ2o0cvSlR3v8vNefvNg
iDIbMNxQiPTq4wz+di2izDh+5Sybfdnm5ulHz/UZ6IAhimkTH3qpbs6VYMyR/yY/
5h7bCHtbJvLGXxgL0bmNUS75rehp7urIx3a9MD5Ln4x0Hfj2xOeUDdWbmKGPiUTc
79Vh1y461sq2gd62YpJAKui/BgM4M2tBuGbYZgtyaHnV0d7p34MNsbrlDfy34R72
ndiSrbyuxF9jxusOjg1A1HW3ym/nzg9EGleSrzJ/512/DA2LaRdPr9dojoFHYEB+
9agmoicWqbKxqM1Z9fn1rsMzgpN8o2lDvv9u7i9uQ/8sXj/yh59D39sBRywwQMbs
+sEPz7CMs+i51P9N9AmL39yfSTe2XRG4a9/n8Ez/nNCCsH3cAXVeDuSMCU2iczm9
gtVvMnzeMw1O6L8+5MR6TbYUAOcWd/ivPeJCPHj0cTJG3FHhfcqDbJPj+HFYddww
QE3EJwSEGwpbWBCTTzYrVIF5JyhC2GfANURVRfRMkEVgwS0SK1Os00CNkzXyErio
hEOroM9mycCvEChEEX0WKMEHNvbDvwLZtkSsr9zmfX/G2kVgqq+fD+WrgHLpnWJ9
TLPrH1y4FpZ9mY5V0Y5lhnmHGZupfmmsRdwmV6Ex0IohXViikphfk2YuODx1Kj1x
aHJuat6nfSD1PRO4FtGTpgehWHp7M+NVot/6GKq2tNhQmDMWXBW8FRApTwh+GOqf
NIpiWOBfzEInTMeSonSbNgProYdhZZI+wF47htbdYNi4FfQ7sJDrttgjXOGqlXhE
Fwz1lUGWFY2MH0qpn0S3Kk/pTweyvQj8rdYwdY1/0SNenkDDPrTK4hSdpMgVDZFV
Qr3PxUUk8Y/YREMZmSxIrBsD0nQHFB7ZFIsmCWFbFVaZ+O9S6b6fzVNFOLxp8xt8
tpuuM5LkQGj4RWcdw1jNIJgM4XZWRgrZAxDHjStoVXGodm62AZYpEpAAlYCrbWE9
gKH91ggCiex6s0zUTu8OpWDjr0pYqF0HdrhA7ksQNc5brzIpIA5AQW8KoIYfZYIW
yFGNU85BrXwc8ILAHhQcOVlcYpErFsleAiShWJOvDALkv+koKxeAebbDAz/qvNGD
UxrEDuBQtgfvDkKuyG+c+zz6YbGEP7duQur87CgQutUcAnxPXtfvXJaU685STuWE
aJlp3IDUYMlFvwoM8Er5yJ3/yvH2ea7OXc12mW3cp6zcO9WfoUo30xsYboF2NlZ2
YiIZqY4uOdK8K23/6oMpvbE/CSZMVFbaeZcHuclMmJoezBLvPrAhdVU5IWv5Ov0i
rPqOBIFt7wV9QHhQD4rBEQ3d6g67zZMiR+FpCE5c7sPVRNJ62VCPH/67kISCNNrZ
Um9Z70GFRvsTlSJTKBnAqcyZpwNJ1GdMRX99/jgSaoVq3swR2qigPB8gQ5UxgafY
HVX2B7h94Ku8AzQKSat9MfRiA4Dwf44/gjvm9A4FWl1XW5s/TostRnj7HY3ZEi3I
t2Knghy0mZq0oqlAjdpMLGiL/MYRmw3s4pmLlttc8hV/lyCT9Evpm0KbGvv7Gfl9
rDIkTZPSzJA41JwxmUqpBaSZoxY9TI5diRq0bknd2yIKsnsq5aGx9RJINR7rtZg/
cWhdvvt+/9f0W+jde3ZXs1rKRztRSc1uOpjdWDoOn5dJ7lK0u2TM4W3aVj0z5Nep
5ATo/X6zKYPOUFH+UgqtZ63V9B2yAOidqw0+NxbUdEEZa96AWYp2QWRaPpNaeBTc
gsZ3tfmW2fqrvq9kwc7DGqYFmrQahr6aobvyabj5fRvwIXX3LqOsdK2eTCDks+Ow
IAonbf2+rrDFQ0d4OZgz5Ens3Ksw5TDZlMWDg/wLQELdW6JgIGoDc5Kx2M0uKL63
rZOQd5SYlVdRqdUNI0WetZpO85bqCdEYbeJqT95krQgWjMTzGa2cV7R1AUJs9p+o
vMLOfT7sgNMLtdgpQmPEr8y3dIM1TkS6OawWx7pNBlxkoaALRb2QwhD8nYspwD5P
iYWcOVHbZBZ/N1frOHizhJ5FDT2FsCs9lEYyT8wMOVP63+gvXeODUEtaxmalszps
NMVtY2C8Cj+YfVzzsO56G4HFfORYt66An41R02M0c5z7wpL9tACECZX3Zq+eqDjZ
y1XbLEqzbZ3IvYr0O4AwPVULWXlKBs5CjsNRDt47/pqKZhD026lBQSm4JioinH1b
P/fxUcs0EPs+w4CnyhZ2wn4mZvuFyvRc3rmk2Jkn2cM=
`pragma protect end_protected
