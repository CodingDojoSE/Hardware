// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
j8SAYXdF/cjX+P289OsRM6d9te0NWiuLf/oEotJASmI1KrKBXRlELkhyRUb1RZn1GP0mEzkaCpA3
Ao6x/YDWDBwgYGAQwSBDlyuJyaDRnNwcd2ERHifzzaz1Uo+kwdxnqurIVBjG8HDLH+Ef69HQ4fkc
Atu9z6Bb0xvln9Yt1NiEvXqtKZixAiyBurQ1pvpS+yD9z1VVmIq24vSZAx40gKd4eWsjlv+s98kY
vHHhrjkJNZzBIGdP1K5auaXDZxZZxF0pkRw/aOIb0HgFbdXyY53fBOP82/ifz+ACnwogrKoxjxss
xIJSklTx4tsz1XyqbODgVJ/Ifsv2H3Z6FnRfFQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
d/hI8B4ab6CPFfc6aQHhQbK4ajCqRlo9BYT+xXeSQLt/lbQbJ0dddUbAsMi9oAHcILheDUAVNq3V
yqg3m+xjwq3TGvcRuuMBbZ0DBFhlMXXTQNJHlb+UEoS5Cf7WtXHH5+T/TEg/PbjVMy3vzf1HCJdN
tcYdXxEGHTs83AJCqEVPzYXsdzSdWjayVPIUOn3RE9+CdAvyobwFcxQEKeVbJauTBcM2yE+bBfGO
sgexGxfNJNd1hEEHXx+fUIvPCzV9uvBHd3rNfD3Zv45Lsi5ShMsRrNB+m3QWqyRlqEe3m45KUbDa
BNLu2dGa4wlri6hrsHIw93OtIDM3WYRvzz3DfTLV4Qfvx7O4LN4fnhcYdjMaqy19OQS0PssCw4yr
cbAiPSy/St+JAWkO7Py0Q17MoyGjrmfynD4HvMAA6UBXYmsrukXCG6ZL4VTjAtOQclSZLUHsKsMW
rMTrAPkA/9yOLsHB+lyCQ6tQPu26i7N6nbkaJARPcDGWzq1QQmJYXZvZlZLvQhGXN5r/9LjbPSl3
B39Mr1xTDc/xHwVvHSWWTX1J20+Y65/TbB9Q1u7dYD7i/0mQd5sysYhtbdv8ussSVZ2ckUJDiVt+
Vpv9xu5jGBJ17Ykbu+t+lZZRMx/ZXOZOpA0L4/nRAj/WlJck2B0z/TCgKIiwxDD7NwR/ayZ4IlaN
8dFsZgRfbvA+om+XgqeliI1t/oSD28Vn8xHMqXPDCz5Iv68o4pO7Q2c6UEGfjTdXEGgYXr8cd2Hy
3fEQXVU+AEnXopKZx1np/T7CNlUPQuLlHjZnCPSIVyiPbEsDFShCTNMgr85xgndbdSwEuoLGv0LP
GvKi6oY+94Ry1UM9wWjj5nOPWKrWMDqe34yQaju0snHGp40oTlvwGcemypWQALZz5Xl3POX/BpHg
CHdmHaUk5bc3fCe+Zj2ZfPNTJEXBvkv7F9EFgNvVjCOj0wWKXWzmYEXQOwTbImJOP6rxKpHxH+Qz
CiCfkNZg/sL/6w7kzpazJWclovMMvS20KRkNOK6+iNyJ85d900f3+Za32hE0nbv5EZHBZvNT1DPu
ooQD6c0e/Sv2nWBUZ23CsU2LPHvuBOfPJaOattJCHBo/faePETqmeD8CBIqiTJ8LUbwBAYPoIH3Z
31593cBWM1/GgDeABcKLsSIxhbts0LCGceaDB4GHg1VjH034rggs1B89KQQAPv+AeYyAB2ZRiRmN
qZEVQsp40CM4BjgamXt+RPvp+mJ6R9zTwAhr7nwqD4XcYelxFs+jlS4wGgo293NkN7SKcEGKsyNo
rKeCf+UflvDn9o+A9Fprzz0jXxSOvkjSJsr+HKnsEV4qxuKkm+7cMLnQ2fLCYfyYmF/gHqCdedc5
D5ROHqItz5+FACzFyQjQln81l23vw/gcfeS5f4PlGVVHShnWHAOhWMaxdfkvrC9p+RrCV7BFqJvg
og0mYmjZs+rZX4JdXZD+LSjdHr/kqxpSSLYpQ4YQxRL6TiCDYs5TrlvU2xpJhg4DelbxZDCv3q9c
iW0zgoP35N+YcVDgFBahs09ne8Zfa8XGj7+yqh0offCqgnn75aEgbfUuSv9to4qxQBWXpUGPuLMK
6OqurX5z+JaxsOVYlacBlCeAH1nOZlnXngs3raMGdkUuzIZTi+VwerIFYSdJquGOArggNUKErJJ0
ZEauxvNxSmWWxxpzDI5rrCsezsHBAt955Wx37WbyFtkURtR8m0hRyH1VTo4f6J+rIz7+BKqtAdZ4
xjVRwKR1JbpxxgixmL0MSUyHdwtWOg1hjk1TrLh2mSR05E/DOwNDs3okSrTbZ3vHGNW0lvgl8yf1
jcdvPbD3pkZVE745MsZvIc/nrUunK5I4u283dS1B0X4WT2B8vjFnEMGsG7MNNcCYSyIcPK0k+U0q
PHpa29/38FozMqrhStCNmoVGix2ruCqOUemAxtb7hpY8hqKuy032cWE0ym5nT1fZ4kdNMJLlKk7o
IrUWm5NgmEYu/R5bd5D+DszpN2Z2/MnlwdR40oITFBIhoGYtcOWywJKiWeg2RqF4mI/zGarqTukx
Wb//RSVbLD8xZPYR8/B+BPhEonlF0Yw+RRSuuHo/anQOiO2dbTOO8b+5uAgYyUL3IcHqU9tspKXL
0vcIpo+W8UsdlZDf4KbumlxYKjV8H99Xy4B8iH9RK2jkTKhRyb9zBWgzfEIwqp7EOx4CQxHHGu6h
OiodAptGcvlzees/dIyDwtwsuIwE/K1agjgTnkq/mw2bTo5U6oGZ8vNV/12gfuG2Mgmp7EweZc88
nvbOp5kgojCs73NpRNdiQeuIEMoIZ5hi9YKKYDUkjE6mEm4q0XHy8nJjjg+baR2BsbjHlx2uSPvr
zxsaFWOFoWOhnvjD+HAhz9TVFu/5hDt9sLcSNzsqJQ2MoTKbCuMweDooBU0U1+U6lrwmZMTqz5Sb
scWmop37QhL1pzsDDZUorHQl/jmmNpdykLbZ0unfAqQC1HcIcNkY/QwwAHSpRNAbWAwujZAl+Knp
RNnFj+6pee2HXK88DUoVa2drHfIvMAGrswu+o/uTRTYMQJxOOuZV7Vl+p/LlHg6p8HhfmA6x8cog
V5CuLcppkBSjSqTb+9PnX3A07HOOqmmWtkUABqjtoAfoHA8BfTbd38QjUefjj/cBhk6ecUGO6pvm
tTerYYqdZknry8gca99QfJeKVfix81EchMg4SBbBtXf4vzWKk5at+6anBQEZypEbrthzVM0l8sme
q3gMqI0WWFyZayhM8pT839qfg6Zez1/TIIXHs0CnTA+PGQwBOk9WbFtKQZMaBPPfcDC5h1QCDLHh
Tk5Fk/MOpyge0lAjOHgCGXH/Zs3o7i6q0YOdhGnXLxuKzw4ZU0+L0S6kACivhakdiJHbj0+HqT0L
V5yE3sS+0Wm5VQxTZg/MUIaVBC8J9h+2Qt4/M3wNmBAP7HZ1dwDvMRiBvKkudS/vO9r1BUBlRBWT
6wK7aEYlKFtSw1KXKtQ7C1XmWB6UoepuoVSxv5SgK/YDZlBUBbtuCfrGF5/5KksWMoI4nVJz1sLs
ykUPYBMYIpBZ8/CESSEb8V7gTdHI4qKlfhNNXQf9ni5gsqubj9vJaaShrUfK17g+yWFucTMDzOgR
70KrHXnRXiv2cq60fx+BEBezmhQdpG3qLjNVNrowvUC8k5a6A+jluraS464Y1Z27L/ZlfdVBVS7/
q6ATaCdtmfTD3l0ltTCqREEK+kgxpCuckAoQlAc9ve62QhSk9MGZgBZ7oDuaSb0flVy5ZKoziCs8
sIyG9oEmI6KU45a6wVTW7Mt9wP11VoJy1pcvokFTcgmAT7sWJnAZPus3Fj6GUcNYYK8eojPjusks
1wDJgZaC44Wrg/VmIpRCOuawSOyLTpxZ+71EtEe+B0I12zgXj6ZsAiSG2gF7mqh/k429wuZ6X9zE
8EuXpNe5k7y2kCiCqlOHOJz8l4zHVkfyhe5cbCQV9KGQEkMc//KKUtyP+H5pz58QfFKEKSzgAQ51
QlNRPOnXyzE9xq2vVFSvVsPM+2LuGkZ15XUupiLbfSz00OHHLd/ooiIP2lcFxz81YRlnhvsAk5Aa
6o8chhNt9HC2uKkGMmOudwrx9GbvWBytJPJG0WvxevNOeka7wquI8GTvt6HrZxhfSnX0eCSc6RSE
OvJPo0+4hlUeWBsjEvju6ohjGxjeEXlMd3G2BBiVYywwkGjql7QRndsWSs7wmJfICjt0O3DPAF1f
/r4iYJyCAgdZx1g10K+MC7+/wY4Srbs/V5nkQx8XoIYhvjhieHF4iDgTAwceL8pjTmpTlRcrJOnO
5VDj/cVhxlqNRUWP8lVdzmqJX1XTnCWKIiTD1B9cfLsqAhm85jp7LCVTP2jJS4SrqAnmeZAy6PxJ
3Zi6wwFqy41IcyYqfYEiDZFOsJN9FGcu8czVxI/boVLOtobqZS7TVUa0c9NT7qJ/1vbKe8KQsQut
hT+I/kUE35+V2+ooUQkfDLEjRTgmxpw7UpajzgY8kj+n90IsdbfIRtuRu2H8hpme322gz1qfFXDk
O7cBeihYRdwSPQ6HJxM+3TwxCb3wYnV7CJmqCuGkD3lvq9sjbyW/q631tkmyY/EU6A3eaASqxvnc
R3fWPpEF6FnUwIu0bIQyfNBuJH5ovHwSmPfEISfqfvOiOGpBjsPFnTykgDdIXPihXV+aHyggSv2I
qB7dT4qN31INGHjfS8WR9tov4bSfoWwAbmnMkyoYFrLl6TWTK437UxyFjnlQxTDmAgD2sn+NdTlM
p1ruhhyS33QinDtzvkIaFxddBc3UvDPmDDSEnT2qGMRMJUnwzH26wjNi9fyQYxpMjq+un/y5WOyl
2WW+k1/CPtP0y0hQDCMElFYUaPSJNKCSqMfLObfeF8TrsSjLDIIf5n4JD6E+fQ5VkaWwCEEQOad0
TcT1S+v3m2Y08SiaFhIvvfNugoskga0uNoQvNiajH4XSTH49UftQBOLBITYiCa4b57SHPa68RYbi
Yyxj8MyPf0Ccj+WqHv4POm7mGIXvOB9GfdZ62GbejN4KUvVXEXHo6L0yzXR2yILg0wppWFfuFSKl
Pwn3dh9iQo/zdCV5MqRHyTaeuqleJS+Yc0EOFK9iJkkhFUlDmVHWtxsYbxCyapgRAhJryxfXaT1r
/bA/V5hi1Gl35AmHMixj/pfSDF9/a7fTpvkBIy3fYrPNbrim20v5aGPurjScpfKSUFIv1AxZNke5
g35e0+Jqdz+FiX8/S2qfhJBizN7o1Pns/Dh5+2qFuzQQTt2ERE2pSp6jyddReWKKZCHu5x+ZkHTt
SCyduOI5C7x5jI+4Zm0HfvNiXwvXRotSla6KcLMMgZ2CtziT79DfOp6qIJwy6LL+E5rxTvf2jhxV
BIsS3dmyk9BoDudduJ4M0OpvUG3qBmhZCdPyYDL+KY/wOWOLfOOE55psDGhLEVQgCoGD39HP6VOO
4ALxMhpBLAVwzwDlb7Ptu2JkC6vIfll3OPLqBzBWHuAKyq1Oqrwp5HebLenaaV7JCY4qM43aRqsb
O0CfUNHUC8AkzZUXxMZQ1XA+PGlB5vgdN31uG72e8OC/lnBnY7q+kb3obM2RSIwwLL2XYThe56la
19tm0xNHV9XOzqWD+UoE4Q57A0bG0c0tBuEvov0Z+Am9eqdf1z3N5sviqIVvUfyNkyJ8pCGBmf4H
CvajWky/ihKlbrIm6OMW6J7ddrpYV3eXdhHH+vD8Vb8LiiKXOc+SHTam8zaIYkSmsIZKnSz+imU3
UqaI+A9B/HZEZFQaJOvMaMn4OebjjUSMZrZHu8DDg1x9CmG8oRu8KJYrWhdszLabNsC9oQZBm+H8
lQ9BJ3BN+tWNjcqLpCtKYSvxK5hjgi7tPdPQ2KIHEQevOJ+m1UQtOn5Nzi3o5aAnEDEGGaYZ6UkO
pi6QCFsxenKsJDRJSK/4/cz+fAcqd2XI/7tVqGfo2IUKwC3RHv1h0Ay0gz+iOPe5ysx4wPIt40V2
86WScL7s1kIfn1CNDqKVCYP/6Bm+VhfCT7yVsHAezz5b9vkkQu3KXGOFK5tlNqFkFKU4GsX02sPR
cpZaJtaAyTUeL2ccFaMQldg3GQBpXbmbFcdkP15zeTvHXSAx77A186SKZxluKlXLIeBBAmvu8Vn+
FSs/KtR9jD5QpEfWBHz0q8SWeoVH5uOlThXtMtKpya57i0+HJ8mLSK2fu7rLiTw/ySehYMTEMbVq
Elz4vAEltoGbUIvcHLhqoua4rQlcSqETDFyI/y7N7+IkPTW2v7vRHQfOjCyxvFjwB8vLX75dV5cY
ZlKESa0LLZLpO/p2bMuiGQOF3GeTbfiis+7/JkBQRv21SxKibaqM2R/p0DsTWRMegOJmhKcCopqp
bTmPheAU9UTWmLpOnLQ+4qERwHgzGO6AJUO1YY3AuBgg5PGijDb8MEO7k5vb18eCwKVNsSM89HDE
in21kgKVUXNUIZQhj+ccAZJOsNLlNe3LUJ/TowU+oFI96IGDM6G8jOPKxvW/nQ09bM4uOKidjNM8
pZVx8joet8UqZn/pg2SXO/HTW2rpbPMAHipU3YSQv7V4q2AmyaaT/wrFZw9ZWHaH0M6V2EANgMz2
/pkD0w+4iLAVi7a+c2IBacTTRmpm7YI7bMmg7A/fpSnlLGWUrOMXele+kKO86Ts5NOfL8WsdYAla
nwzN0I+2nFe6ZTqZh+bQzlVkqHEZm+SDPESE48DfpsH2KoloT4dHtESzeKW+nZcNQu+GuTpBzK/S
ZaFzJ6o5YFzdB5ni+2fLDIGecYJ3QZp06BYruzzRFyT4vYru0+3vsBGUdQMiWldVsTebvLManhWl
pudjCry5CGab0fbYlZ4rj/7jGaYovfRBS/qfXieYQoUb2eZe+ZfSXXbtjA4J4KpU0ZoSOjEPRjvM
PG+UDK5hrbr5PrkbzBrq7nl47jlaJB1Cu0ZjMcRkczS3XNa7qJyIym7SvcXlwhEjSYgbj0Rclafp
ybBUFzrdGe3YFrNcaiNiU3j4xYxdQNQoG3/vzRgY/7e9gv6WBq5UNRWbmJKQIGUNn0bk3Ye8mjb5
FX3mDx3+Wz1ISOLRZVWqOS+7MHS5Zg+hjJY0rZEfZkdlZti8A5jvTZ7ZdKpJAn7pIvo2dVjrGsuX
YU2P2OaguXUb2vfX8kUV/IUf+vtdwIDvC8yHg/0TwIXR/djK1kpEmW7SebxkU1mQrgVm/ItRclhA
jGyXbj8pEj2G4rz1bBAv+GzAbFWpmpajWjoY1vMBTz9ZruuJ7x0VfXCSwjSSYrY77ra5tOzKMNah
ORQsht5uv/nqMbT1WXio6YIt6pmEq7AG4lARX0F367RZhCFfclGyX4J1H8EnK4qe/iX5ZjKxBvDK
XdgJqsAh4PTN4qCtUr57oPkXPcVUQ1nBZeQc+2I0pmi8SrOKpa9M3i10nj0gPYouCEB90GRAriMV
sNm/fcI7hsFckLg/aQXBOxCPyWrBbFWlR5jTUb+XKpVsHjXlY0o7hpT9Z6a/PxP27BBuxeud0/Kq
fNOOnjJzDU2EhHWBnOMkYLmYFSPZ+45BnBv+hGPgkIqMWe3KAKADcjDgblDce8brI/hM2X9sqmk9
Z34Rz+zFB7PMlJ9R09IWe53u+/hD5p2J7Nsn1aMRT3GNOzjM6anukKd7nXkxbJsf0Naek0DMaEHA
9pMO52/AAkZ6NdmwK1u5GVX9PeFnX8k9s3XyA/1nfzgemt9peTy7zXHjNfFhLDbgxZ4Chq7Lyocj
/gObBvQHPKGoWygbbPsl2dNXglvQUaldjR3kmcOqF0FwgvXpbIeKajQyULjMOnpynPNn5WDnFPqs
/EShRHNQU3ieUCYrJXFkR7CcblW9A7ZzXpSJil3OHzjOW/v/Hv3e/9H1cb/lu7Wy00OqMzVBCcTe
UB6jmfh7bJNNvifwjNSVVVjRRWYMjqfVDN9O5UMqvCKVl5zWnJmWU/V7Fqw7jzJx5PYnv5uZWsAM
pxOT9E4j+cajTOIhhr1ZCRS+CGyI6RFlAgxUuDohjgvHwhGD5lGf9l/E8P6F1US19JzRRnUdrCfl
+3uJUcmV2NCpBF8J+TkW1CENamEYmFQ/S7OEJoIPpBe4a6n0nIzIKb8d68XylXATfC17JbGwCAO0
MRbOiooXs/o4kyQHqpNxAVL6WtuKCv2mtp8g8CDIiKvdeZTGZHMCEMS7daFIGR0QRYl1Bo5sRlKc
kPAMiiSMTROTCMPyJHzYjjXHme6wKRq512IAa3aZpG+2L43hNXwfaqWbnwN3h4ce5Ex5IwU12ZIw
Grs5kXb/nMnzM8SJiuxQbdG/k65JUNlERWbN/iRY4BLcurMYbdlZacfqYpeB6az7lxvNnMKg2rgZ
c20HpNEwo9+fonaemK7stKePTyL6+Ed3C2UwMgmppRfNw9ZdwukiiMF5jc00sLUEi08mc64V1aZ5
P7wYBrXlFq7ny9phci3HK/RnT/OlbXVeWyCWR3tS2GD3ewk+uBNsWYSL25KN5q59E8eQvH5X3ycJ
XqHyvxpfCbrDrKrCmxvNTSrtT88TBcWvkjsfFTU5iQpelSs690V961Xq/nDVD7uKkKkp93ewEbqm
MXjH8Zh69JXyIFz33tWxotWCDYUPOo6xkMq1jsbgTfWTvVLYpJ3Ad0oj9dWzhr0TnNkzyG2L0hxJ
4LbqQTEuceh9Tvdq3Sn22x3K48RILj54GaRhPVdk77h/Ad+YxhNZovgiMd410Y0WaLAuL6ORsyph
axvUl7L2t3JicJSz7qDvXPnGwcpScrCBbjldvmOpMUKJUO+oe0WM4EyZh4OGzwCZY+dBp6yXeLk9
95tBaHji1ZjUfDrk6a8d65ZM99lHpjsq2a841OtQpuOfwwq4gjBqddw00ojzr4viJXE0itj893ZN
EmLHYRGxTvykvx1ZzqfV7E0iDvnr7kaF4vHVDaUk+7C57yRswDiJl7Xv5hIbwZ6bVyQt+YcG1Eck
ax089XAvlg7TComeAqTADhy7XyVx0YWCL3Er4aImXq3JUj0zKc72kIbBde3iSNjtJ3xdUyY9ucPq
3Yxwkn5+jzj1w70oquhQ2NTKw2ebN4kTnxx9+dJAw9X4weT3Dk7+Au0003cvZnjQBHs7wjAW+3yO
P96WvOuGf4ZW0JgtOjYTUgHgPtcrBsw1QaE9jid/RjcZ/yB/7cg4VhCo4XB+oY6f4HQuEuH7/HB7
hZ7jVGRemv6+Xl4f7kjCwU67y/LQr5fedelQ1OG0k6j+KrrOAj+0KsK4EP4zZK4IJ948FwVwC//9
xN8YTtiWTvXAORYmG3ACRF8CkMj37TKE578FqUIN2aMS5SQlcAlL6oRxJ72j8dn/xyC5/AeY4fal
wXmh0XArst1o0nCbhCvbxlKlbWsBaBxBBulSsFiO9r1Ls8tNH2waFBlR1kmB+KiHPHIbUjfBmanw
ZJTxJVLpagV7HNJYNBX0xfTCWjRdG3e72dBvlSjlF0wB3QX9QfimOwCm2MjPCCt44IwenbPixrGD
lsInxmWUaMiKEfYArhcpvB1VmUBEFik+kNZ8vlSQV2BVIhLOYv+jnbjez9Lt4GOf3zxmFaFEGlOc
eWamFNuSgualUNQpJD0RZHjFuUvgALkSHIJqehdOpFZ7FHw5ID97n39RcRwFJR6mJUcWIsWLBf1s
5mVUk3yScz9/VuJEw0ecY8Ej4BZBwz2ydbep6ZwP3ACnAlzqqaCwRuMMxeaX1uKO72S0v7gFSo2j
u77nYx2tt8mppVlR0MAqKZrC0doJid5yxPVx69MsTJl3HqkDbNuQPKRf6Y/5DuN8m2s4u5yQT3ty
vxHpiDRLBd801Ja200tDlvme6lXaCpfqmSkolcAcc7g2WfOKHZoGBunIeBC5T50m38ubaxG9InSV
bZ5W8LfEjK/lyOzMpTjaqIV5vAnV6frgTeFTttjzXiHjVaZDAMGy6enBifD+l/BYrbthilNV+p2G
nAIUgA4VLZ/pq5iEhfGoQ3ZuAf5E7HkHdo6xDt7Z/LSaeL2i6vRKg9LUMfX3X29ZE2rlolWa5icE
7/sUKlwTXoB/tMlg3/KEWAAEOk2dMIgzu+mpVZRa7iHUS87cZk6ttxN0pkOTl2QYHoV4zMLOX2DU
mdJ7sucJP23zPlrgmwDVLiGSuvnjHMu9nFpN9kMFJfK1abyPG41XB4x94DIZND30rOQ30AN6jyG0
PVH39FnuIW1isRX9PUnXhdEXIUkBhVcHc3pMWKpDhZRZ5A6lVzvL67jWFHyZTSgCp4H1xtS8nYRj
KqsrpOCjgZt4fuBgdNdJ4gumRYu6oUxln4qbDxBX/ojQbL6dNaols9/mG1tbyoht8/Mtrrx5KxPf
mTNd83CxAZh7en+kS1+7RiiybOoEpmNoRlsE0iwBGlwxti5Z31+cPCys/5WNG+fRNc+FOugs/ydA
8HNZoY/sPE6AMRyx9H5en/Ub0RaC+n1WfvcSU+DPwukwbrQTeAiNoMc55FFmWXmW255MmVLWIuzg
bw/J34SIWIL4V6oaYy7LJ4UiLYEoK9Wn2gdBdgob3oMf6ZGjcPvpzC/V32Cw+aLBXdw1xqZkVIDL
h9P/OX8R7Rh6BcEq+KF9RSXjJEPlBVj/skdqDevex118LyM8qmwc+I8iuvgHyDXkmHunzo6EHj5r
r5zjdK2r0Cul3Ms5xbAjQTGgRkdmR5qnxTnrdvm1iQ1zMLti7P9fATyhaGp38tErki1iqa6RhlPd
0ShPE/TRD/L1ZA4CApKdmMqEr/WdzuooaC3kvdXRiGqqYQAqe/k8J48iE4l/ID7+yeW2wsiLv713
L9oKKRtEI60epRBzmp9yRe7GncUMdXM1gY7IwaOoTqt/jn9Kc37nujTx2Me/W9ziZAyTTbvdNcAS
VSawDgtbospxBmPCvY6Xk1eY2Swu0U6e9JYDY7jynhjXZseL2eX0t8PmB+1p5+LdurGNcT27npVy
0xURZqASjNOEuAVPIFXW3DG+8Mz+W6udmXd/tzsIuzS+hUgkPr7e/nd2TmCn8Cb88KhOFpyfME7T
BirpRdJCuKfvcCsytuZ1qQgQH9OsucbuBqC/GscflOYHZqOqKyYxfmK4uipy5ZCSRERXPbK9GNyW
VrBSgofNkpRgDWzS7mus3abGvZdgssKZJnYtxcQ7GhIu7gRYKJxeIQRGETRbn3GyCnZREFbedZRg
cIKyVapaw41KK+EDnb6YCAGK+7VfVMuyqt36XuPYdWbSzx/hlVqmBfIoFa+XYwosSMv/0uqLBLMj
YkoKflFgp+lRc70CMYQBS4J+6ifV1j2Sr5VyOUOorX90MeULYj1yHa70ZvuigCuehIojl6lNRTve
v41oI1z2WRuPnUqMgEZBAxSyFkvdClUO+zqhKv6BfSuiuzFSr5JgUkJIPrntnwdqAeHIbPn4Zwn1
q4eWzwzboothOVfbciCxbUutguoVZYosaGflApfbq3vVNJhIDdg7hcqBhrtyysT6Q/4XTRhBl4iy
+zPx1VN5njWo7i1Q2y3duCSbNDbbSf3P5CsGx/lvvXvpZU97yhhBb7jrn3Nj16Q0uX+eFQghZhDP
nLdm4a4qdz4rJLNWfAEmFfRuHntGCZ9VReuavAaaC1l+9j5puW/PHffcbH5YQ2XO1KaUtswUQBKK
XWgADi4VeVfoP8bQf/Q3+6qQxQY1n5aStdtWJP+CfwV1AuC+QVaK97Ux+k4QJ1Ptu7Jvnzcd7rL0
5muvQY7ZkAv05rY/QgfzuSi8UtxhSBPe7EdP7JauLrTmJInELVHQBPbVuM1mEQ877Evs3cVanYmz
WAdrrARBZi7AMzbRMZPN8Prhd1NDmAqGL9bjD8ZX1DyV/zR5cBfGxE/g4Dqg/lJ/K3pzawSxsdWD
AwqV+VaBP08QCd2UysxWGUR+xUQyvydjewAkXzti1Rkde+QL2xOpp4MM2FOYJP9BlGFjI5Lp1HlI
10MsiwjtV9BU/nzUUZaSe9rueYz/A73qLqQbr72gCish3P2KhEqN8WsDvrIVpLdfveTmh8asvsk1
IN1Cnck0z+cVSB12pSiy6OSK5BZYd30tNCeTr9phdBKz/WC4trM/VOqB7z3W7TZzVpEe90S1fsR/
6SaOCtsmyE4dYBM1to4Fmm7037r4F5HbN2I1qjxRm9Ft5rmpaZyiul+28sYbVjuXRWOvasvucJcD
EzJnoPvlz1K7qvEIvXAeLSEJkDQWJH9zaSL7hhHH5GVRtjYhsGQOxjVTgR5PrppbBpXSrWhntFcz
L2YG8m1ULiZ2XcHXrNBnv1bXG3XL5DtfR6MYJOCftlTsf4x34PnjkXXOax5WFRhEdIwICtZX3Euy
JbJiJQR4hnoPGSbRuoYzMoOQjmCPOIdpNjO3jRwrcD1P5vWTNiBIFAomgHuDcg5/mahZJpWtN8WF
/IfQBIkGfhWRehOvaEdYFD3Bcv4dpPBNsCk6Rh4y5jzMNA0ZEcu51YTqaJO+sDx+cevMHp3pIvFX
wqkUR1mhejF/qjdo+gkqGVzmod0Ko5jnxB4GMiMYuBLNSH2foA5/ikZBXoSqlz1/l8AWDDf35sdm
CEbQc3mohKMwVY2gtrLibeJUnZbFh0O4ArWkElE+PLtTSuD1cVWz0AOv51WHwvueP4J4NWM9/bag
HeFfduWMa9fWDQJ6Hb/Ub6lXXPEQqsGAm4LF7XODY5JWfzCdI8AQeWS0CZJnLm3v0RGJoy9egyqY
GmV2oQTenLt0qzakt7J9XLaxLked/VAkvQKXijlRW3Gv+ZPqK5aTMKbDqgtR+R87DLpQiA55QURv
FPXhdS/gTrsI/65dhM6MfA/rtSuiuNkjhDmaob8JHwLPJUFh7cbSRDeDqy020P33zJBLnemEA28K
J4twMYFS+sbdpa8p2tfpgjXKSPH6lzr1KkuP+lSOMlo3DUzuphQH3Oxv1IcmaU7bueKgB4ifLxB6
j+i1u5xsq1/XV3BEKTyydzew4E7F+tLkr5Li3bGIZk1ZDTULC2no6HJeUavnWp5ZxeZ7e5LTr18A
rWhJ+xMCLyKVaUVLamg7H8usn8JCGCEMv/XRDXKcwKc2yklPGIWR7O1Uk2v4xrQs31KHJd+Hkcy9
ni1gxeLjC1yLeSrkmzo6Ij1lc4sXsOVAABJqWCnzjiycgcgOUT7NCrRUJ402D1v5K/auw7fT1Qsh
M5Y5FGNfvrnRF42jRWGcWo643uGPtlEGj5Rf0GTNUDIohVXD6nVNya4Mh8OTTPPxCcEHWB9kmV2+
CsmXRNP9M7b8rs4gU7P7B5HVwA/c5Gf9o/8iDrtIVqaEfxc+4KiIrOh7tVBhX7wUhtbFRmPsZqDK
sFppqGKvo9b+nG5GNl5YfLf0zQiUi3wi95cDtar7AZkcp80bJrO7sY2l9LZan+832/EOGz8RdBFa
MpveIN0AiBwAqGyfCpLk6KhBY3n5uIC2lmVdm59A4zWQaBqUsW9ueIuuA6oQEro4ucDroP2xztqa
+jywViE9KYOfo5lgCO+jwQa/D6jsrJchpXwMmPvtbqv9Jz6ta10YOEbF9UGyyQkVKJnjyoQKRtLJ
IMr/6m7DL9FNlycebl3jRrWRJer7yWr0H3r9Gw1QuxHII7Mo0Rq0L/ETk4xRyGFpCI8KVS9oLC08
CmM335oevssRRMTZcbWFLyEu2HC9H9QheFLq8Aylqk1W1yuDdb2mwlfPz/s9/aT/lHtQNmQZvuMp
Rc3u6rbRcP/XEkESsrcGKw+2eAXtWr3OrfBV+a9XQ4I843n4t0ebm5d3eV2XHwTr41kpGn16w/fP
e7gbR9nVy94ECPYslNHPr2l6XZZ2CPOoz9zsej1JoDjMYawRtcRc4GVY0aXmyZekGj2f6YCIVZbc
XjgpLSBmgykzHFpSRlyCi4DF5rHcsjyBZc/JGcyQ56VM4ibN8HpsQzhc5HsG2x4405YEYgEAmm31
mCKIWqmbiDJyKh1ywZHO933Vncq92Z6DBTAM25k5MromIQFsg3F3wscl2bz3dujkC/CRSEtmipA6
3qL/xHJRuGaez69r0qV6wl+6XzUIYN6DkyN1ceL52wjkFAzZDXkOKRY+j/h2YXeuc53Z2kfEKvMh
0zkUSLRk3KSxUTQ+kTvVH2vV/jk3fcLTxdadrImSMBJ6HpHHGLSjN59G7+gGsx0daprRfqvXmCzs
PKcm3ZTwrqdWgHvdhSrYzdUSIf68GZC6eXUG0g+prXhUuvp78MY2H6hez4ZIb67neM7Vi8wQ+++W
wxEW7hgJJR8kGhWMRzilOhejMMQRpwMoiYiwRI5hQBUAcGgqe+2T2BC/P0hPdRkGrO+yIx4eTKwe
63K68jMfgVNXnEb71iNGuLkRYE4/PiTdWsZZ6TDvsCpF2rvk5peZqYPwzojg7WdKVuNyCIwfZujF
hEn88KElRcSs/LHT+4ruCOiBj1nfzrWT/rBiIw7S7AHs2yiN2u7Kxp6ga8fTz1lRF3C+sAVadB7t
9/qjWaYll9MPuVfmobhG1ovdRbweBcEDQVprSlRCrONOdhEdCZ22pi1peaVOI16iCQa+26Uj8P5l
mPXv9rAfzhbmi8ETYhgQ/JIB0Wbu92Ym3wIN/yqfctlrJsLon57gQ6IkTTUyhVA3Kkgb9rvuB1es
HbEuv1jACCPDJr0MbO+ZfUN7jp0tOKA4p5kMJKY0Ge5Tq4hMIwzRznGi8nRhYtQaHllMgLeEmHLd
Ld1J+JH36bIEViPwBXmOjeeXKK1uCJvPr28GUYJXfgGMU2azrluMtg0J5ZcKB97hJU+1fIFYdHdX
W3Mw1BARpCCTaoex+7vnUF1v0bRKO9Rhx2esmdXzRgDm3UhOkWcvqSXn9RRATPvlM7jjSVP2ml+8
mG9kAUTGQ768P9GOt4Ew24BShtuLkBGwCFE/DEQwK2rVSoD2R62cMIdL4XMWSVzMTuto9dOKVoid
gqP8NJRBbdqIlcCFnnRIPWeMkrcvcOjNnKwe0vG7UItLSxYukOCq9w+BRuRgRxZrXpYlhgXqzwfF
UzrOQcsvzLZtAo6oyzzJbhxAfpW54CzaAhG9XW7wCG+P1OZaPDIqvjnxltSv3JbHB1PL7zjorcmc
+dvOF3MAu/F+1eXnz4kK2d6T1AFiaZHbiB+tZ6unrYGMX1la1zVsW73HYG36W8QuxfTLY1f0bG8l
Z9W17InOqQrPaXBQTbsE8AQggXNT7HHy2g9qusCyYZqNRsnz90CwwMWQQSPH0duypaTHOtNVHCGR
9ZqRm59MK797udj0fwWWo8DIfGTP94f/lpI3uWZw5NwVSI/F6Hbu4wSx7jQa6JhdCWoBsjUkG+WQ
hcXixvmKImqyFbt+T74T+/3RECuV/XPyUXTnAjPuBkEGJFRSfhk0tmoVTmebZB8uTn3MVp07JSLw
GYgPdV+qNu8CwBsVp6C1WIqu9USF7W5Xh6RN+JuW/1WHF8WqPYT6FvSQ6MuDEFcucpbPkTZ6swAw
sjH0MbdOJRNucpp4hDZ6e5MRzgqoOEjtdawXH2rNQ1gpRoy+YNbBinBYXNExRyeiLu1MFYupfPeW
3P4nyMlWt6l9AvvteSuRSfo3xrHEWDSarZCuMeQ86V79zDh/jfbycceTbvKUy2i8unl+pnJRAfxg
s69zGG/gqShH05V5z96IRmEeNpGWB3aAdmsPtvlLUAktz+2Dg4dZglD/Mf9PAa067vT7c+ZRLK0j
EkqVlPtWt2+yTGBCDiDphrqM43G1scljRW67BjwRolSWV2yET9REQAJbI4fJyej5cygoMUZV21pA
70ygJc14X4hyCVdCUAN5AzbtlHBDIbxywnIk7D8psNpAGPWJTb67Vw+2F0MuogjZSeFt2i1N0lRN
qpqE0qNwi2zPVf7PuDO8PYqbhKPbesILgtrj7xVmiaxa08XfJBstRLaf7+aufuoHZ2stgE38af43
1Zk3hd9P/jtqtsQgtXj+GlvyxpCa0qmAwnQacUOrvffTuyHg4a1ZR6rbo/qkc5xBRHRziQ2z9WEg
U3acbFqDEbFMpITVz/HSLkD4WTlJHKI7Lk7uzzh0i0I5+kY0617JBqMUHbMHKXwtFL1acd/IUiTd
XnT1yjIt8AhqO9J+wuERRXsgcASZVFR9Bj3NLXtFXs4dzVBdSeipv6tIZu+e9RzPtJCsYuVZ+XRh
kxROa4pbCxVHOJISoC4ldi8yG8QYSVd0zgl5IZHsru4QOdoXdjFaICs0neU6RBDtxpUppAAfU11x
g4v2iC2Kk7CEgs4T0y90ccbxcA/zqBiVBElSPWqfOAywahPlwHah4tLSIhH06YGELvNVQrAeWgqf
lYsfouFyY26ZqosqYkU5Abg9mXlHeAwfcEzZcVb37O7o2cOJdcPdumOHyGHtp+puQuw68v8gINTN
4ShmPovgARl/8cm2KcGtHXTRduKbeuwAEgyhNdFbJEegICtZMMaXpKHYrJSQTsv+J9atKFPXZBds
OZpjboC3GhTXVM1+I+pN8jngULy9xu1cZtWA2oLKNIJPcaMlt0msStv7fhY0c55ws0tlF11e5lyv
O+Bkc2NW4eugSKEtiRwcAFaz+Yp7PhxoSeLyI2xBWWxVHIvajCZdHuS4sBdZcehxvQ8qojDs4aVI
itW+Q6BupRwtUfIdhlcnY/77XBrcwFiPisicxKDEdJoms56SOTAZrnVnIXnqNstfF8+fhgKujGqP
NqO4Slp3NroJJIrpD4abVovdn5IRDXRjmRuUfUteQdDVmpZTeCed6zslzTnwYFHvuIkvKnyyCZBC
PaT9hZChyUTnTklrmt0Z5yshmRtRSxySKiSMHitGjQKFCQDwhqcN2I9jiF/EHQ6N/gFuZfgwGTZn
KfN1PSXMNCkk7xF4EAC4pKK/hZM1TlbiOuRtFhYd+6/gYC10sLq26aAugu6dEpk+ALmnEG/UUhp2
ONbJSTNz93kLnYHEfABAKlcQfrJlchcCkwbCNGTVriMOeC6nvAkWXrwEWaYWXS4b7tcvOA3+hyvy
I6s/GlVFpSA72GEv+o7LCRn2TQHWvQVou7h9JlRU1YwTeHyp4HSu/a5IhlYzLb1KQgE178KV/WsV
lhL7NHz/Mb9/GIfSuf9HZ90p+DFFBcZlIfMQTRE9Q0xMDKOxAeZSAQmlkcp4L3QZzRhvNoNoqdd7
sg559cmOcu2v7uGQ/nqBseU6LyHrcr6tCIoonv28s43ePjYEqJW4N/7LNqNpeQg7FJJeHmFMAeib
VReuhUpggbQ3EkmSzy0a6D/EYkPF5NmoL+SQRZC052YfWW+EYTxFX65Rpxe3Ys95jDA6HFWmSET6
b90MMwCrAUfMF+mHxSIMLwH+ALI3wltLJm1rn9xBiSTY8iGfhZseqfS0Cb5XlEPGZ24q/KnGeNPC
M6WqbMBBWU+rjDgQSacfl4cN6sdiAFpNiAeYl9AW/aSAVITirALfPD5r1uH4pUkcPMTfOCTRFIbI
8PB2roS0AEjQBRMMpvjOC1UOzbuxDXE+uzzfu4F7WoT5gNXWIETqA56Hzr9PZ2989Rk3CfJJH5J3
pLBHcvUqp0t3Uq6pDzDWfuZwGzXlzyRnzhwBmsQIn2aHGbFKT0YytrdN3SXsvcMZSmYP5/ZXWwIJ
yrskYes6j+/pgM5Y+yrqlBxo7hHL1PYxkMz6vG7WyjMRQ+6qFeMB+pg967oi1pxmh8uso1zhZNEm
NUm+M0JI5LXl1O68qlHqp8tZrUmCh86JJCEsWR9ufs6KjpaJUr3bM1ct5GI4dIsB853TPH0kUnC1
wXuEY6ahF8jbty7Mki8YUq+R2rZ0zm2Ahs1pPsJ8FrvfousACGwinjnYloZMULwWqQaHb02veB4T
dOojC5hqa8uGux1KdGtvf4DelvW82M0OPi33RMzgcBVghj5B1tuUamaX6wwppj98n82QvNpR/lXZ
P/f0WXSTJXRi+BKL3tj4Xe0tsXtdm+dEvhnA3lrvcpO4x/Ugt/j7jAHBs9QOgnJk09j05ZZkQRWY
32sM+Y+P2cFWf2dae47EhvOwCJqwBGjJjNDM0l4aDIRwKAmepdBr3Ym0nvbdxAZIQCHpDiy2oors
YZr+sDbodExLTpewWD9UV58PqplykmB9E5o6eU5JxA1ZI0HlfZb5TfEEu5JmoAyl7W3XMNjNq0qN
0V5K7O3Gxutge1aDC4yoS/l5D8oyLXn1SyL6lswoE92JVxVugaBKaPed9uk7kJUyCw7/sleMGVPF
VGByRZvdhO4v7fib+mei5jTmfGWneOwhpdWzbbrqdb3/1cUhPFhWlyJsQ9Jj2P+YRALQ0sRDuR/D
8RGaOyqR/K8lL+BT6ltKb3y+YT7s71s8XwVZg8j1IRbfev56SdIVyJ7DWmmS9bho+un71tadXjTN
tCFagHRkp0QUA575uWtoiZc62f6k5BjzsxYzl/14LbM6E00bmiUhhbzFEP2vON6MGc2/lgEIo2/f
s89Y9EDs8JfaYWUcHdaEMn4yQJHManKUPscFz8szwpBeBPS2FJdMnWl5Jfqg5E+vROuFp1rk7z/r
nZYGHQmqO/iGVI2U6qQgBL+VN0xxvQJmq2XIE6kVsc0qJErsLmPmtXEIlWx/bMBFfuDla30AfYBm
tqsfRZHT4ZD6jJcozmjrM7fk2Lp9co8ZtZ4THFh6IajPDGGwuR8/qkCN8wgPRKxrAZcPNc8wRjmM
rOYOefvum24yM/CjrGyh/odvJqDXY1jPE4jtSdk6CGQURSzDAdcMGTSyIqUqfEuEeCJnaxcJmEkc
U1obALOXxIqrDuOgE1zr02Xd6OnksmA62ZorzXLZx5PakweJrKIGKfYkOPEea34ctMKn+2DDuBO3
51wDPmlSGboRCjdFaEDhVpL4T15gJ4FCWik12Hco7YGZjdmxt1OX/p0Gnc2pr34npWI438UEnzTh
R31zxFR7t3UV3PauR46QBOsEXCT+oDp6LzeUmxrSRE+uNosM1f3skxENlYgm/vNAGkkSQi2AhUcm
gnUB8Dhe6e0fuXPCCY2ClHInMRJ54F/clILbUrEnDJvyw6yTq5AJXAStLL+aPynkXtd8o+RwF1Fv
ChIUKw/Yb9HJjlU3lmJsvDcAIgzaipnmzdo24+E0Nww1JPCtbzVfAyuIJzRhrKVgytgIz7nOxSX2
s37RQ6Skkw9batZFHVd+dcXo7uc0+EQwrMvVZJ8aEpanbr5jPw591WAsNI+77xDUB5PTRzATqxIM
HMx/M1zE/xeh7dbBrXgZFdYEzBVZdG1NawgzkP8X7VUUnWu59L62ujEDOyaEK1BbHf72xLQILgFU
Zw7iUXQD+BCL4LTe6s5vFNzFLEK9KrUGmPAaNqNaPtc3ImA8xb9d9Tg/nirRdj5jN64nUqxj76FM
6FcEDmht5nThmApQ8clkq27tRRJxqdQSHVAGrlASFnljaC19riDg7BsYWCg8x0BqBtckt1jOJCon
p7YrE/6WLoRl9JN9JH/fdtiDvhHJjAlyc8gChExJHSFiZ0cL/ABoG1sviuG1Ge9UWx7rV3U0IlfK
VqXhZUf3ajmOugn1eK2JSK96bkXCy6XEECc1QJH43hgZ82gHghQosaBv+0A7iEERmIi1ckRVM+mv
/a38Q/Dx2hivZAQ52JL4H5fq7pLZcGhIa6CZnCHdw9jYdV9AnYvo/rwV5VRnB7XYEve6eTenCB1N
IMw8y06b8T3Ohnybk9vnGV8zAezNSuLQ0jrGEyihuXi50tFcnVC+uu4xVQPNmspn7H27JHFLVRrm
R9IT45E/d+YjtY6fbahFEf8kfLxmqgPi+ptgwQpmMHPC9Huf08uFztRpSXw/cD8F/8cPtLYkpr1G
F31ijE1EC/hnN0n+nbLq4Dm634CZHylLljEZRO6tGTEGUpTKHanap2W65rD4N3NA0am7eyJiSgrv
fEmD/UOKvq44SdcAyP/2+OtNKOahfSnY0ru4PmgSVSzmKxnUXCdXE+lqhsLK2lCSHLIoG571rHuE
TAlCZ5XCEnbqHf9F0/UiVm3ayZhvi3tp4Wmqy6Z0elYmbO9XowL4xbqiRbL1TEYsJVP3Uj0ZM9XE
yIGHFyGv8hH0NNLbo34S4xwKzhrmO6UJ2x+MTXhrQ2T82A8BrvNkZCMxwjzK4kkS7rbTN/7fyVyQ
iLT8F3Ol69AnOjc8FY5feEI13nwo2insksdHdpaCtsPRhQ+A/6aLVLZCB+na0wIV8ptORyrHdrIH
pHADdUWgl7JFVYU8j938hIhdEWqb8ggoEVwIAVTTkc6xZivnxEfq0acD2DFsAWFoKkmvKk7o4XIz
sTGDKNgThAXxrJ6V/TuTWIZ3zOetty3Rxa/eOGhJmcASE0ka1/3U+x9s7bUwQSX/vcrSEhQoGT1f
yo3gUPxNoo+QsQrg5fgx+VDNF/dBAUW4NJ5S4+1K9XaC+C2KVA4BTlqVhEEoVJ0QADCrJA2Hp1cy
8u1V88QRiSzU8XaSN6c9Xnc/DW5HNFZjkdeKi2pFVly28Z35sfqq2Q3BKcKjy9Ttz9g7uHBim+/V
VhvVgw64jMCy7cLfqKW5w2pVNFERn6Oq8kaNvZEJ9Ouyca670IDOBTkN3HS8AMYM0gvv4TYksa30
p34rADYs+wame+F0JeFZP20E56YnpV5pIExXYuSx4CEV1rnbHVzhE6+DwF0o9DRnBzKtWN28nHAU
nHn8irgxJbkU+b2YZOe04p/IQd/7GXHUVtjL6UbntTJFYgNJ57ujViKo4Myiz6qMghek/NR7C4Sn
+CZfpu0AiBDGeVee4BfKelKwPhbQl5Q6ymRNC4E0FZknQTgwLiph6R1QPAW20kS2wKLKmnflBYcu
eCNBWLrU0e9Ge/0W0mGdpQMhC5lAeDafEUJmKaY/g9twRmy/K+4Y1OEsvv3EZVslYf/Xg15DoH8T
QEORRdca/4fnBhGD1hUIRpivTt0F68Yz60ISweybAS5q/LKuEOrUDFcDEeZdee/LT85Yx4KpnWV5
EOX3VsTy39F+UHWwbASIVvMCVCdy31P3Dj4oVVvL8JcUm2LO1H+Dh2s8JaQl+T1BUVgjiUh/Vm0G
m1+ZoEDSs6qUm8MKtA9YH8YhWCC004s7xmhrq5Zm9qe6fv1iBbRoIbLENl8FUsOQ4qT0eC8q8F0P
bHDvBQ8ct8JKDB4/fYBcpTi3iICdzAst5MDoOptc7a6Lx1+ImWBDSXu953F+WCvf3s0A/leHjt6S
eF6JdFxff5cLyT31GtIeKcJTnT5LRaSlwy286Nv4Y4WA/Ec9S7RansTFPyT43pA1o7daplZjIaXb
2Q9BvP5J6ruymN+7Zkf5UmgeZ4jm8b1JjyiQoiNrbqwJ87aSY0m0MR2T3rKtYSyDY8YXhtr7EMN/
EiHYvEDU7s2imtHl5VEqzKvPeHt/xAgPRTmH1Q6twvimbeO9K2Wko/x6xhwIWJZubO1KhsVnrVQQ
KvqyAbuM8fw38HRpFdb0Vo6KTj05y7rzZawZ9wroSTetG5XM1H7eP+d965DLa9ZDSr+W12sjpalg
9icJZvkoZLNzpFlVLgch6I3a3jZ58y1w82KvinPJlhRcmAnj+FksZfoGslZqBJh7I2z2tI2mAcHF
IGq71aoe/yfZVHLY0v5ikgKV72LPPi8Ay5WKdoGdcsN22Plh5inb0NwwA3bMCHsb808JK8BVcafc
lAX/NeftwWrdaBU5nOE1pfCKHawQ2UvG4LdAtTWu4jpd4j0yQlC9lOPXjy3tqnRSfAHTNxd0OcLA
5LGAJ1UTyJJxcn91YfzAyNyUoO6XaCWyrxXBCSjUpoGWM6eOqaiCqdlBP6n8LP1z0wgGsCsyrE71
gGVIVP9agk70Rw9YQczI31RI+Yjgp4EewdC24x80ZlBiZuup0/VJ1luW6Nb+I46Hb8cb9PJ7ynhg
svoRrBJV6VtqeRUMLBeaEDjc8sf4PkX///qBJqvB3inEY4HejteFakYoE88/p3a3hUJdx/umXVnj
8juoP7ofsT/CEwobjEqY66KCip814ua9j/l9CnPfj9R/uHD+q7qPa4uxRVw0yT+AkZbCXhcArEMj
vPjeNnveF79vb9vBDNfkMn0Qz8RaR1w0ZejINMWdYtHaIPvu2ln1LLoGIiDisHU2pO0Hg93tZbH4
eHowaKnb6HH0B7HTwuvAgBF35N5Fukpx2ooMDh0We9oyLFwXGWhLgitkbSZCwbqnvNGS5MqV3Awd
aaSH1hI9C9ARkm4jLNF35o58dvaJtCHmbBE7X3IMssJQ2vwFBvGu9+6UUlumOgLSxeOu283wYX52
j8rw6OAdB6U/vKd8OQULXMuZ/Lsvb1tFBEyQqohRUqSyzBwuK33xCnrttSA3MWTAz7xgZmCCY+mR
6BqdKNfiLI1nkIrysxBRh38l+wydc+uajhvXdHnPjnEUS7sa56FqN9Gs98nA3uw1i5JuiaA7xVdl
kkHKdrFrj88km1GFw8gCFm+f98urDi+GG23kBJ/sUTuxUfs7Gb66hbNbKNknxq8Z3lO4pFPwkObL
RhvQYzqnbf44pgY+DvlRNytLnDOTpxrsfc4KqFpqUKb+9qfQ0F7+OT+mpqxjWDzQv79PUNAvKi5g
t+oxSBSnpZu2MyBgpXNpX0Nzh6GCZu3mkAwYfvSWbec3xIJ8xgVw8Tk+K/bbgjCeGHlqR/Ya2OKz
M/nTXux0fIeakJsKRmP5IIZcanT0XrPKRBK3MXs1mu7XBBp/+SBSXctaxo5RDeHGO39r/P2I8cO6
POmfjebY3ct9D4T4U2hhy//UdaFkichJjzywdh6OVB94YM1QSS+K2KbY2JiZGuY2Y0Dmydy387vZ
ITNIcnpyUUcNhFNwzvwtq9AbVEaB6FGB+sYMN+lUg9YXLVJLPQfnAM2Djce47CL4RPvEuYxSEIvL
dKn92MfpaAUwzRkUsZnOxFwFVxhhOOxjOV7vQ5u42KLhVybMvzPGaBKGKTM3WpB1pejUNQQrd7lE
tyaObIdJ3Ej+ofsW1QGTIPGzuOHtbAMnwtrc+WwNLlzCYB41uFtgu8ZrFkW6LVPS2pQ15wYKF4Q5
vz9j4W08YFf/Z8pciluZhBXB0inzcIdnUETKQ8jy9GfdcQcA/34+J0UxO1PdH++9bYHhc15ECzgf
cRBjtTye57SAW95mOD8ir1/ekVdukm7TDMyUSlr1qR12AgoalIL1u2BDgHAmhxcb0pz4ciaJfC9U
zgD9NyQyBuDr9pYLs4roeNksupIsIVnLrKeaNTQjFFj73mZRWq+3725+PKIirBIsnaLbaWN1+rHe
/Yo+1ul/E5Ksi+Zg2SIviBymxdljYTq9keY2+R8sG/kaj6z+eb3gOtVIj4gBCPPzZtbMwPFHfrtR
xCYFb1ynKM/gkZhwMYVyqpTcdXqypGMMYHf5VIERv7VzIEK5pnekzoLm1HSC9NfEA8n6hjL09RUN
W5DEoR051SYHYRYExcsW3l0KnP8Z0KH5gEQH6HdOBQnD9WZC0VWAbWYbmaWNiYGA7H+twmDBmW6j
+8j5z7nj5aShhLrvY2eVhVzD8+ziYTEYOMflE2fgkcOzdCWWXWgWVyn2XTpYmmF+feHrP7ifk3gM
Bpt5iVzbrsaZrxabiPDGPeDzFTjI3E3nWI3n72n3CVRktAQGA2toWDhjhAccw44Tlr5IVYdLJONz
QF+Ew4UqUN6RX5m4pK0YiBApUXaWGEnQkBkOWtONrMOxhWeaYrQ8Jl2nboigXe4/OS9rv/GsKLpy
VEVFqjECDWyrNnVJ+xrx2ECmd/t2eSQYIcwMcfPDZwsQp+jlv0SXKslgUlMRvU0z3kRlsGzeTGnA
owGFxFRitI/WaIYo+RLIZPJwP/1pkbbKUbQmUURKWcw8j7/YfRomVF8bbs9tSiLDkMPX4jNd+u7t
+2aUX6/MfHP0QB8H5alNAuu5sw5xnliYRwp4Acw8ztIgapYA9DWVfNPbC1LfOiCqFqGplLj1bhkX
2YRxkEY8ZNRGaTCAGhowvEW2aB7rjzcE4B8ZfvkElHr7lk/dCKFafx734a2u3nWMx+FVec01FAK/
KDdI27b19Qw9EbpRWjwxXYN/RlQ2pqvw+a5X+iBTgjPmnv88XlWpVWJeIKa3opoNdH45hJ8dOf1t
GOGOQVFc/vkA0meI0Q8XdnVr9kSsGguI07LcdRSMVXpxYYrTUnGMwtrUUKmbG0pYDw2T/17Rn03B
vIlCkyILo4d8ovqIPt0gc40OdLU42rvjNK2YELDQ0CLbf5lktatBRgkMMcEvIc3QcziCW5GzGtw9
XO80nbDw/+ZI+dLR8oYqpVC7xwH2DWEAr3joqukTtdQxXl7aM3TDpUMAI1TdNjOhBZp7R+mnjYsC
OExZM+/ZBXfIK+PVMyuIQ2z0ZriUAfi3WsOvFIeLSucRFMyTjwnjYUnJshPRJ4EfFmalkzcB9I8y
Q2odopzzne88NA1pwuW963guJl42XzPBXfqHiG9Hc33CibsX1k/sTVB6aORONKheC7aJFAqeLMgN
vYeB++OIxa4JhFqveFtHBlK0HmqNKs0WbuxfAtlj4NiUlkxiPr+MRzL3RDmHV4Tgv9eJAwxZHUjy
E92A2umMTQjQEEJMUIYf5wG4IaENMm5cu1PmUuPjwqwhkNorjHBvd0w0w6YisOrR4kr1JuhrhrTO
LP8d5SLQ5sMETLI5wq1ECIRJHFf8fLU1gkxWxoMzD71KuwwCrBXPqQJog8ovAbSTlvIZLexNWmGc
t6MHmcWofAmajeDFkw3+6S8aBjBx1pR30DAOGMPO/Ui5Sy0235BzzkeDTTKlU3TMPNNsCSOgKzxn
SPp0iyvqLdGp1/m07QMK71zIOtZQQAN8bZxWteHEljJb1x+SDeOEPPHhsHUndQ144iPmkircPHzG
GFQcgCYGqBGACwySjrJJimzfz5+VXyX+B5epNCnS8XFM4U/nDF7IZANleZit35BsA++k0ptXydyn
eHQ+fH9/SHKnckYwWqTdrSJTJ1ffq5hWbAZXTBCEHdiQRCtQuE1FzjHr4ztX66Pva9JdGd6igkNA
rXjm2r+a7GfWYM9ABF/dzjkE477e8Cu6oLpOXkmnIFUsovje0+fa0GCjI7XY9vSsctsd5/W8BhcI
78WIYBiYsMGP+thPVgEGc2dub6QvOHFKP2gGwGIG/ldJn0+wgmg3BAZmLep1hC0tXKn85k11NXmk
CZIWo2KY1FGpjDrhmZWUvN/VVo83VNVGpBEzK7J5EfDNV4vtp2oEKQ1jUMRBBRtL0G4jZClroh9a
VdeyKrkmLCFzurZQPZvlolekrhpO3jKKe65monYaypy32TXiQ9nrJ4zEl5tkNBUAYQVD2mBs+V/J
b1ahownbJi9ZUkwV72dgW93Bm8pPPQYloHMJpf8J5UUFtBGt7/n118dhYiWy8uh/l4YJxuuf1h/q
3aF10cvOG7N90HjejXbNMTMVavNQobTPcGNlUYyTnbQ28ABfKmB4TWfwn+vfEc9VTPYJIafbQsoE
ML4fTNwArZGmwZucm13djIlGwudQtCYmpKUd4vvP4Lxi9ekx3/eyeddwCe9O9sHfFpSWpYA/D2Sb
MfTAaN131KkauvtEt9Aue64leI6jdlp3tz/Vzg8ri/iylip8u8zQSGjyLhhEFrnNaGEJAT2yQyuA
iM4h0Wg0AFITjcst6nsCRVJr2Xzwa5BGttJRbLNzzWF7Bqi+rBrMN4MbvMs6FvdvPa1vIJyqMZHM
xDHgcK8Mt3W69FfHLUdL8q9KyBy7m9dwE15RjSMfqDrt5rp3WpSPVYIMYSNOst1u88Q+XSHDlkAC
y3t31bjiMRoUu+IfatWRlQMMN/g1h/YyeSRbRoWAhDt3tuCs9MNOensGTVq0wgUQg5Kmvt9uo3Zl
5uikHwVWHVw9BBRqKnxawZ291SuuZ6++0n2lhkLBaPPhCWLw7LArdxf4fX1bTF0jHUn4RCNyJpTq
eKvUEs0AbkOzgx4FYyFD+E5fIp20bVCqHZ26aic95q7NELkWxd0X7weqdBIqMpv7dpVP22Wol3sk
nxMbEzi+Ufx9WsceWk12tRzFRNPFvtuM+Vdfp3tYZ/k7ij6hjPQZU/uJsY7ipl/eViviFmJVxIzC
/cb8wk50i3JGhwQzB1MZWQ+kG851Nk1vRk6hO6zFvl9FtOTXKvzjJszSblQAbPIMFemDyOrRXTNs
9pnyR7Hfyspsv79qMDW1CX/jhKc5/RQUtucTEsmGvK7NKCdDFw7zUxlLb7i0fScdTVdG0z3Hj246
D0V1VtBI220JdFdeOywRLxFrLS/vzpdfZTkGfQDX7nX/M/GmVV28FFU0ktgbPGnVl4/1OlCmchxh
oD/IXL15r9oLA9vJkXRMc+obOnSyqEppTDJMPgwePHupmfSdxjGWASVnJ+KIE2+c7Qqw+U+uGE7Y
UvvoElAa1I4csJ78ZWzk2uhqp3HNzCIw3/W+2jQ6sopWh1LlVNhrzvwz+8B4XV7te4xhguU55S9p
lJ0brE8yrIvFUxyKKubp5jTfnmMDhsuA3ClEk7rHI9/7o9gCII1xNvvqZ5+x/dgNJ/bDVVqyQR5/
BJi7V581w8yVjbDAaBlS/jbNR42g2WjjGtanTDk3o5v3BuSaYwJZUIJmdUv29HSz1xsVNJCiR9tt
iU2vBlTt5ccn2l2n+lu2j8mqoQzyIfE3nilQxbQTyD0gNsqbtiHK0CaBudyhLhDAisvR/oGxbOcZ
AbKNsbeZQpPdtrVee8hz5Z+zBvP2KhVOmnLostKg9zqtYD5RQzMQN0VLaz9hB9NZgLSdlLwkvs72
h5+NueE2iECXfuSUwv2BY8qHO4pOrdohEbP5XRFP7wG45lcRETXRi+pNc8L75k0CnLAeEFW/S+ae
mb0g9ZnufeYeHNeSxUqi0CIz7KQBKol0UiNU9/WUQmKiRxX81FesWWLjL0Th/7MLmUMCR+XLLDNP
PlRPVQILhvv54g7MYlv/dEjJKifa+XBNYRquchL5fYfQo/txgJcQshVpxd4Mr74WEXiyXFKZU8+A
JZgTEtawW5n8y6NPQ/LQWIGY+iw0T7aqTjmoLT1v+QtSQpVL6owS5kHwsZfS15ZDWk6TBaC7adSF
nrSoV3c+VKB0qMxZbS98Mff2xCFxepEWv8OAm2bNU2A87cVuQXrH/gAKTp5CT5+gGk7JPWmSgTsI
ZcwY6xF/vS9NapvRMdU79gyann4SzrdZlCx4kVm4fMaxIhChRnaSlSU+DUbCJvEXFunNKI28wmr/
GpD+cKDEv+TYRZGcgdncZ0/Jnez7djmsT57HYx54CQ/qaH4j8MgJz5axbr+vAUAj6k6MvhJqNWki
fiSelZ6OyS2YvCijhnh7ulTNoVCo12r8mdYNVxwrTHCTePGAFnJTa643JmcOUfsd6NOSbXQH17nB
0TSXg+tkYmaE77HqmrlqJkdVAIZHNDt3BgaIlenCq/H98YkVAQdoCLRZZzqVzmdvAhJwEEuK9EBh
vAHMVmmErIFNZHx94t2H6D1y3BjPmIjX8AlLhViEykGj1nuPwWOw1dlcQi+CLOl5SgXvd66PfeFF
7WYgTdoy9zk4ttqtLILuNwpCDUU8QiZ+jtEcQuzeU9uzyM3A/WKBwuz576CN3q97H42nhMLsAgUC
Yi+e6KjboVBhxqFUpv43+OPD6ipYtH5BOQ2T0OjM3hYtuqyXhYjR/E1gIkOWbHQK2Dx4Sefv2Lrh
m+3Uf3AC/7R9nvxeIf86C/MLULDsJcp37CfEKQGH5TtwVPdD1PrgUYihP/GWZd0qAsTLWqyLCAgx
0LGREkOXv70WrorTqWwhqHrNX0J6WRsEe/YvV6K1cSucTBYTloaKwei2mwsj7lQ+5VfE
`pragma protect end_protected
