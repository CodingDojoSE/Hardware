// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H(CN0HTGH\Y1EPQ:&53K+:__FP_"N6L8O5*GR,'##-3'[4]!FK:.$-P  
HX;O^AF+<Q/0Q["FP"#T$-K/L V++(B0_%74#J4MKM6\R:&=:>'C*MP  
HD?%R"NE ("@#&9GCKR2S+;\?:K-4/"A%T0PU77,Q?PT["7HDL"#3,@  
H>M#W_K92X%^'+?>-1J)^0H,UDP=(#)&$:FC(%G!XD7$GU]1^5KL3>@  
HJ4A\VW@0C;W /)4-S^20SLG[W';Z.HGV&=0LGYWI61D/N?>83?(/#0  
`pragma protect encoding=(enctype="uuencode",bytes=9152        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@22>0<4.-Q))T"?D4*^)CXEO@9!UZOMJ0C:B.W:'<=%( 
@IPXC+M";G%!P2 G!SX/X"Q8EU44>*7V"[];&K%YCO-D 
@\M&\;*J@/AWIB=4@QKK> $8R1C*[[*;Y 1SU82!GS9D 
@00%Q!";\:<=R)_#> 4(_-P*NX ZK\ E3E!:% 0]AD9H 
@$F1Y*D5QXP'"BYW<VEWS$$^,8\W7'0RKIX60._ZA7VX 
@-6/^4W<>22NP=^7+94<8)J-G &XO=2 ];@P)Y<)H$I, 
@7OJ"WA=@MB123O4Y;KA3%SH:/0.R)&?WN'O%J#7+ !@ 
@>NNZ+/,J5ID(0&+HOS,D>C3>3\!-59YX[5$U?$@["7\ 
@RIU>:WX?&M_,FJH_&.+^&YT+J^-7E??._/+ZMFA"6A\ 
@*M^>N7E(H/6-;K^%@*QC;XGQ7,GGMX/.W6SM+.M][WT 
@R+!X\1C*PVRVJ5S"2'S,T10#\I?%[K-, 4<J3]UAL T 
@W7U4(.-C:7PD\<&Q),5[K1YN)11P'^B ;9O0:O>4J"T 
@#[S74#0@7"6-WH<SN=U9R17J^ZPG,N;Q8L>U6T'WTI$ 
@09"&3&-,"Q$/&<L(YK+MD%EEL\S7)N,+3X)=[XGI03  
@J<34=1T:V$YNV#(KGTYR\&[VNFOF%A&.]#%#35(3Y&  
@M'@_\. B2KD59QA#0UN4)R&U/J:]%$RN6AE!L*Q0N;@ 
@;(3A2_)3I_9]2G-6%KCRJWC-6=T[-]%;VM\*S/$E/U( 
@KD4$S8L39F?(0(+3'&4EDMCN4[8V0[C:2JK2H28UCY\ 
@HRIBK1=KZ D<8QTXL+;B?XH,OJG742^UMTAG /2@[1  
@H7_DP7/_'VME+Z6DW9-* E1ZA*.GQJ VUCYF(+)J09H 
@0E5'YV-JV/[&D$=@8])0\L1Y9S/Q2727.+PUEI Z0<0 
@^X>E<S;AV>11$\@(YG0@YL),L;9M4JXPELWSA?7XOEH 
@:!U(H._^Z';)CSQQ7B1I?DS5V!!(@,$^WBBC?4]67U, 
@=C0* 8Z]N>O)<:,-N@H4N*ND>'!L5(S5CNUW0 JPCDX 
@"N/1E/1K)L/3%W-LB[F?>VHQ_OM4>(E*M<UFP/3M'+@ 
@T7F@P;5\;H&+!^.Q+RZ:HG#!4\(F]E$B(KE^<#=/4G@ 
@E:8@FVG[1DP]*M(@0)Z\A9-Z74AWOI[YL^]< "CUU?, 
@17[H&2]N-#".!;4PH&WH>9P[+%SE O//WMF6?B0=-NL 
@1#+U_Q?DQ&?JL&+YV?C39A4K#WMCVZX^RFRHI=+@EU< 
@O</\6)HSK:E1<+NP7TP#81^I$&!/W6&%_+RZ/19NUH( 
@=_!'2HO0Y+C51RP+O>*:23NSE(2%872(T51CJ.9]XMD 
@??4B[]Q--Q.<[89+D9NK-\&J_+7-:7:WTWS)BI;.!DP 
@2TZ$'A ($0FAB/#=NHCRB[=3^YFHF*;I(YT^>*.J/_L 
@DM/J(D&BM]-(H_!QP;_NM!XP*5VLSLPWE^G,^&Y7'Q4 
@.>Y#1C[$=;%>XA'/RE3C4TU:U> [/E=QK^KZ%02=>Q@ 
@6&H&G>3Y=TU]LN'^@[B1S>*3%4JD'EE[=S:,1P4T2^@ 
@X[^V:DZ\3_3:$LPZ<\,9^]3%]5APF#UO'.L'XE%U470 
@YB-TA>,:-'NY<UX0DB73#?PFX=M3[%3/QMU"B%4=(*T 
@[!K*U!#:%#D"$T+</KT' UP>$5!FBCYD+]76TJ!(H@P 
@Q@9$*-@J(\R.*+*8R-#?Q2D"8V;R ]OAEM-%#M_H=<D 
@[,&E:6>&8*A471C%)V7S*<5*:BL;N!_WL?8,8<EIT1D 
@60#+]]0=)0H%<2(I'SZ7>EH1.5/.>81K2@:)"HK 'I4 
@V@0PN?-N8HZ"LTM7M-X;!W3M,0H?CS'JU^FK]U9].+@ 
@(R+:0$\LHNU<>$8A>RAK\A0HDFF(OF1-6SN>!!E6]Q4 
@,KO+W-^1@C@$/K&)S=YP<1:5HB%4:3"Z'@[)<#?671\ 
@4.@R%>(?F3\*CP/T:?PF%6V. C-]?G+Y+U\[1!7%T*4 
@N"2<EBOWINAKC@LP EJFE 2X^ 62&Q8@<<-X>SV1\^4 
@I/LFW($#OOMC^6FV&9*!7M2I=B74_VY%@RL$E*CMVHT 
@.7FNU91FNZT]W<<J#XS+0E#Q,EFKQN[T_X5 =..87$  
@/F(YM]IN;H(4CDZV\*I&O1!X>E='XWQ"A>R+O];9M=X 
@@4D)#27:L]"HI85W/\<2 >9.&H&^IW^\TV?^7Q3%*   
@(K)?#4;PB3$1XC.URCEHK9?M"?,4/$^'C ]V"3/)K8P 
@0&K>-+O=BEGBSFF0@5:E@>T=B4FC2EB#C5S\9PYL.W@ 
@(GQ&JSW0&B:='EM_N!&*2#15VV\+\8Q>5"^46P*"2%T 
@H6SI##V&1T;ZMYJSR,2%G* *J/3:2L>Z=:L#^@)Y7Z$ 
@A>))<H?RR4S!=F?:#CFS62O_8H]B8C#6Y=-[,%X^(9P 
@+?D:8]_"WP(03:0/M:)SO;)L$<[58J@^_A&C78GMJD\ 
@\X^;7"I?Y($S3'[-O./U+.XZ!-E /@O:A)K[-U_>P8D 
@0PQ&G']"U*/5(9?8E[W[=>7EH/\,>\,#/GS803CEM:0 
@"T-PY?KLBLC37,0\0Y?VI +G..P.(<OAO!U?M6-Q/$H 
@CE%64XR[C*WPI:JVQ&@5:?]^4FE6Q_DG""A(^@-.\2\ 
@JUTX=_OI7ND,X_0 GG2@K/,E/RZFE=L-[]$.GQ G[XD 
@ RX#FE#LW,RC0&&90=TN<A>>:WN2Z=%_H6"1N.W,XKT 
@CD/*57*KM!\6_&4MO^0F1/I]'D?<8)'Q6]\6L&7:J?, 
@U5V!C^HX*^,<)C%ME<U<5Z&.&[,03@_Q[YTEW-LX,U0 
@7ID%\K-5_KXE:LGU*_\IF>$$@MULO[2W]OH@!(AS[+@ 
@AO%9WK_EGO;5;K5>VH^AZ[SN!#=#V"ACZ)3/Z6,9S3T 
@6%0*^'>*$4F#105'",-%2YP]&F/?B>@_FSH)LZN@3D8 
@CD7RWVC">VXA)M:7>$J5GK\ ]!=>9Q_YK04$."$:'B4 
@K[E$I/\#XI[%1T?WKT\>#O&-4_8[H#7(6PKS#?O46,, 
@Z' OT<E]A?:]F^^C\@#;'ZS,2' \JW=\LUV*S"NM]!T 
@VLYS_97O0(MS-&I\$X;I3Y,6\X'"67[BNU XWM@KD<\ 
@+7'\U@V-1H5F>UQ(82;\GGT_15^>;)C?7+XV4VE#MW\ 
@(7OO%9I)6$1$057-D_MJL*R"^Q+?6,IBP4D9)$5OS-L 
@335Q.-'#F+)JG[5T92EF?@5[RA6!6V-9430U@WI$>DL 
@=!')PF,Z.-B51UK!BT?S=,74-RA%?+Q*NSNXW)L.OBD 
@>C9Y!N;9FG &AOB#7)GN#]=(LI.1IX)9L!0E0&;S,<L 
@XF41V;- +HD7'P".BAGUILJ/?2Y+3]ZI<NMN\LDBNA\ 
@*O8C_$C%GU8T: OU?8!3N<*I'$6JO(H6S[75Y)O03\4 
@:./H(#"GY0F'LLH[\@P/)N=.4;;1>TTEX08V<8XELMP 
@#P;L=9G^/EG,27F/"BCKU-M.!M4M"O\16-Y558.<E&X 
@III]D+S).Q(96]YRR(8C3X\U6\OB\=-I\/$!3EP]Z,@ 
@E<[7YK)(/<8'WYUJW&TUC2OXTU ;'RR])BQ'MB0/M.L 
@[C@2S^14A>Z&)NP^^48(X4.(-U_^DO'K5,>9NV]4Z[< 
@5#0.N1:#$:FJ_9PYV#<L[N_S6 3)K,]WW[+5G/\#V'P 
@"]#*FALG6M^3LXZP^ JZ,AT"K9'Q2+L/HK.>@><Q4LT 
@RK YYE$A6=%]K5Q5C5;5*\:<YO,N:9+.15G39#2->0H 
@<&I&\$*WT#@-YW^2VP3BZLIJ!5Y@ZOGFVXZTL=H*6<8 
@(Y1EG2[SEO-C2.1_2R9)B&%F,>_SK8VP\<5!]GY$8@D 
@C(I+QT\,BGDG=7E5;^"31OC\&#5W00JR29>]K*4>I50 
@&@E+>D"GF=!BS+8V3W"H#H"LY@3?\"D]0$HHI.V^<WT 
@GWWV;2ESS388%"2 ON4-SF_>EW)T5; #J=@A<^/\"U\ 
@X_W9_;4#+>5B89X(7 /OO''J)F.0:;Z66BCX%LZ)0_8 
@/(V &!I XQ45Q$T\""LU\.;"32VV$^8BA#BQ#9"4%;T 
@.CJ,#-GY_QH4U(N?"A62=W:<P3TJ.IV6+([R0*-F<!( 
@=K45HO,;39]\DJX*)ZY_.DM6AL:%I_9;TPH8 A<KL#@ 
@6PNS+SX5\9Y\;9CKZ>@\[T9 UQS3\PV."927LYU#6HL 
@SN?3==&*]R.5-*EG.JS]@. XY%B^"5\QZ7KY@/(,7Y  
@S@'O EOY/DM#:;U?TQ;+S2+U$B#Z!K[QH5RUY1YS)N, 
@*P6U< 0=1F*F 6@6CWE#LCR/^6FGY!F]8],CB9$^='\ 
@0[?.+B8E+F"O8XZ@\G;I/EXG4CYA=5C9:$7$/9^##_H 
@<#L97MO#SDB@X GMYOTOX\/092?='J^(VM]> *"N]U  
@P1IL ^N>7W&3H/_P7VF=@07?"^G[7*/0_8RS&:%AJZ, 
@S_/HZ]O(N..XG$Z';_A. >NN'<HK4$W+6^B(:45JEQ4 
@/ZV:D&XW-VPI&4&:G8QW X)<)G3*?D-TX"[#]A-5Z]  
@R9$6##%WH?;#E G;N]M'IDNG%,3NSX'\KW:0GVPKY]L 
@5?-U47,SRY5MY:(R9HD]4O*C.#;,";^B:SU18AO^65  
@C[ %$&4A@&3I_6(KUM]:XX*'GY(7--1N8D6!NS&C7SP 
@=>,)K)$I$IVS?%[_$$-Y:\&.6]@,*3<(!$M+FM&6E]T 
@U7@&)G/"HV6,,#C@@1?PW!C*>97N5*8=+K$*A=+3/S\ 
@-Z!%];9W>@O*^(K2.:,T"*T/][PRN6KP' \)0R;4#8H 
@'[(HV'@MM%3*TJ\?\[/D.240>QB]>+8$D;*(Z2,^@-T 
@+W,E%3VWODJ?<_I5!ASGU8)?G_?A_]KHE4<"B]UO<KL 
@*V:-#^^NH]<4Q8;MC.8_TZ)B%]Z+-C,#\DX.&Z44$.X 
@5L;5I)5A)\@_K*6FG-;MT[1NUB+IC$1$L<#2A=\*>Y$ 
@9$JK4]\_ZRHUW$,J+5$HA3Z%'1]8H,"AR\)O^T1-"?T 
@5-A!9.Q$+\FX(MEK*!58KW SJB:Z:5^G/F..'&U' 7X 
@L?%!@I,'ICA"3D[+C?_EKXEK $I>246T924^X4$;V$P 
@8,;*_8Q\W<L<$> )'K$ZNX982G]W&8T513XI>F**JXX 
@,PD]W7RMZ_);4"H[Y#8-"7\8UNJ:[>QUB=#V6UYJ5\L 
@Q"U.O_!D!^(BD636]9CJM9@;9J/<DH(B<M)%?+";?'8 
@=83!?J=JFP@1'O_Z552G*?2("-IIUGE$%_K\5.)L\!\ 
@60;,0J'80QAJQ2=>Y1;Y4/=M JCW1&(:&PRZV^I'%X@ 
@S?^UKH VO+8C,,D^#*O</U&6$>Q[7B! UXE!,,HO]_< 
@RL,J> LQVY9L+\5O7PQMM05;$%7$,IPU7+7/Q-_VO?, 
@V=N[%I8EX-WYL>M5E85*ES.#=4E=YRH0>N]^QVV5Z\@ 
@/IN@ 1X5TYWSWP.]^7E]>@AL2SCUYPJ(K<"0+(=4[ < 
@+K?A:6K^*1X\R@10P4EWFXHP74@[.S$P#R^ER+PAL7P 
@@*''HZ=CE_A4YXH"8W=>!3&V Q60+68:-$FAY3:*?[P 
@FE'4-T0%61RQS*<MD8/19;DD;O(3DJ@\LCAU1)RL'ML 
@,+[_%Y\A?YO ,5#P/;__Z:E?0[72BO-@KSS8UIFUK<< 
@X6_)QVE%!>?LIR(5EI\%VX+)I\;MQ>29,M%8#C'F;%@ 
@R01F"X:O(#&!)8C51:2F5$AL"2/U*L6EVM9I+,IT.-X 
@ *&3[8W?)(X;9)]0"[#^KP+_\/I<91L!OZ+L4B#='JD 
@8DS#;'6Q&C-(,0C)X ]M"+@8J\H)LUKQ#-RPA15O'X< 
@5!5B(I!#;?Q(NGF;NB:8D^I' *$M(JZM;4"1CN-^I_H 
@+1BY$6:42=HMM?8[J"\MPQU3$.5)J>FCJ?FCTC-B!U@ 
@7,+QS&#R?6 I5LW(JB00I"77&SA^7P,0'QJ,P[7EA&H 
@(V0$>(DIP F]TF[3U')+G%"S_-D1SK>/A C526P_RDT 
@3B^^:.07/[VT@Y8FN8L8\%*L#ICJ"L)4UB:F<22"<O0 
@%*%E3#7J_Q3RQ\N+2O+&8Z:-@3_:7$H/#PJ_#,V2 &< 
@U[$'/$+'J7Z 8 NCK2QY[87D@3O+N4KM8]CV ]@>OU0 
@&1B:1QA5RG)?*^S#E5$#6B=,?FV-5^G^'Q"N?%.>3R4 
@ SC23[9?8<R$9ZC\4&5$MAX9.G6I#<8IM](O^Z12X6X 
@;=4HX>*T#^LO_#PP$E7EPBG^SY"K= K,*G]@S*WL0*4 
@73;9C?@EJ?EA$@7W+?$H.$E2#=A*S/6K@FPNRLC$X"D 
@.JA\+BZ'"J8Z91_GP5L,!],YK??&:1#BDO,/9-,^:S4 
@N1^B^6UM.](;/0('\XT@F;H!6HJ(')PC*[QOBL9O-HT 
@0#XTJ\1YY,;('J312K&YO?\0@YBY*R=?J9Y@I;.F<AT 
@0C(?9/1<7NJG^2@,68?84B]G#<@H'FI#ACFL;X<7_I$ 
@P!<#%>2DCN*B1##(C@O6-O[<%47^TQ'\Z&L;REW>#UH 
@@N[.83E?P+1.;,S;RR?$48>APAB<_?PX!2<:VI;B'6P 
@) M$ZR\GL+5L2;7=)E>@;8X9R5#G2= ^E&3S BI&3 < 
@[>IOL6D-(MU3:[Q&H7:YL6?^>JNRM.*N'55(ZB?HB#@ 
@G,%%V=R_@(!*Q1E^$]3H/X9+0LUH/-%G4((F57.WX,0 
@&U&[]C4.^=E92D:,JYRSFQDK8L#X@528-.FY>4OX!A@ 
@HD6\ L%723<&  @&%H*P 7@;0%:1YGIQCFXJ\1Z7;O( 
@YNHL%6P?_^Q&(<+;'&]_-650\R5;9X"7!TH=3N:";2L 
@J])E(F4I<3W. K69*0N,X:Y-OD)RC3)")Y<TE>BB ^< 
@FHIZ-QB19%A;7/A7"R=?"@4>Y?1\)8C8BM<ZIO%[K#, 
@$;N/G;U>8B)TR4 SP.Z/%<(> <DU$I2_',# 6J<V$8( 
@VH.JA/3&FK[UP@9RH!43Z-W<C_Q/*B&#.+UC*A<D[ P 
@?9<!K2.5^A*U$I@\;,"S W\9:/U.4F*2!K%S5"._ ;  
@$%D<(WMU&)[-.O\. KM1D(OO1'J-VUI7E!1,S+Z0J>@ 
@V9C;X5[O35]NOAP6+H^4S6#QH]6?ENY" QVK@ZZRZBH 
@R+0>NW2B*&-6%:!H^?Y$_L=[&2>4_4 9XA'\?\: :J( 
@7V,BDL_75_P@41!J>C,2A\9GOUK+L,K^9X4(!XSKG*  
@1!/J:KA(9AWY"0/W5;/="LV$9A\K7J69J-@6T((N0O8 
@J7V><1>=RF]Z_G:];7_\0K1+^C1-BC-TC=WHYE"YOO  
@R/0\RTV8&46(N5J=(LD!^HH5SJ92<UD43_=%[-@C6]4 
@V$,N*"DGS&V4(@/ BE ((6+[CS<P.'@NHTQ 2>.S$,\ 
@XQ KJ\MN13+=E2#O70R^4PT&.4QR7BCRN%%_LFY&B,P 
@I&O\JY]&)8X4=[Z"HA%^.SZJRCCQ")U'NZ $&J#OVM@ 
@K>:8%<QU&I+NT*:BAGOB(0&]MUIJ\V-S]<3%]3!HCTH 
@(L<A.;C*VK)'#K=<1_^]TG^#HF+8,W'X7?KOL;YYX"H 
@V.!G)/F9RC:J[IP.6";(#B\K;T]T[EP?$-F+D</LJV$ 
@9\8OHS+ .<J7KM&'=*L(XA))2K3T;0?>,D20FV,TY;  
@FU_XXF=R(_61:0,J,D%4 M0,QO-W8I$ W*UOTF([;,, 
@4CLL'D68*Q7QH:*])Z?N1^@YGDQ]M#E\A\B5O)GR4YL 
@[0AB[ND"[V^>OK!FDKU0'E*0E$W6-'ZYB_T@^00P\OL 
@I9_\ PDEDU=OLBK5[V.;^B05[&-^I$^)?K\NLD4$#NX 
@,]\TR(2=.X:0ORIF%?/VWRS>GE>K-Z@%"D#V2'5& ;( 
@Q^E(9A?97&VH=O6YG5$(ZY+.EBRS4ANTL'/F;K0,&]\ 
@A'M-7_9#NB*16G(V,.,C=A1FL 9MK(^%6N@H%BT"!50 
@,$&>@NVVZ^*27^XUZ&Q82=>1S)5O)[B@(4[SZU--YZP 
@0JD9F0*,@D"?]:WK&)JT$;:4G<,0>[B;TP*[5GJ4 QL 
@YGH+W8JH4I#:032<863@CG.IRV9Q?/Q.&8\F]O DB/D 
@)7#QQ,Z!SLJF!!(&HK^F9B55>W38@)^U)P'0'DSXH%( 
@VKNKD0P1,JJC(< ]]V%+.L^D.D3A,T=%VF 7[H7QVL  
@FC!I5FG;9@#D\(,."U*?Q">3"1W*6F%%=XJ#MOBO@)4 
@<+K:BGYK7TE_<TW>)G3D/EXD!FE&;1Y6?BX_)?VC_<@ 
@*I 9>=97JOR.XV::0A'P-LA;,RWF]08<A <$#N$=@64 
@F"T^TSB5C1O6\,S+1W^B1NFU4FWV/E?[DP;X742XC;T 
@PJ/M_'$XM;AIZ?BO5!W?:Z^(2> $\ 0HNA.5\#0(L/4 
@*?BV1^E#A@-%+$$Z!X+J/'DV\L:S$B7[#1M5QF%,M"0 
@+N1_"4Y"F('O'YMCU&3*)1,#K9;!#IL-88H0N@KS.J$ 
@;4ES]4DZF.DV=_K.B';Z"9AW^&6&]\D-3A!P:OXQ:P0 
@J(<;[SO9S J/%1DL0S3Y1?82EKH*3/%4X9 RMN3(L!4 
@ _/T<V>D#REB]*8L68!U+("IU;DS1%Z)^&%B)L8N"4D 
@!B><S8#'AM54#G^?1IY?4UZH6K]Z56)6^0! 3O*Z=LL 
@5A5V>@Q6\=MW"*=)1NP7_BP0 0O  CE/GO&!S2([)1$ 
@&38P+<\GU^7?$WAX&3V^JO%9MOPFTC2=!..B2ZZQ&K< 
@)=BYV;Y(AQ/3]3;V<W#*\S!O^K\W=X1[XY3-2.90U.D 
@5W[YY)L4LAVRFA\R)NKG()5AN^N,U747+=-$[(;"NHH 
@4(;V(;EZ-5TEQ'O-47UQ+-B*GK_H!K>>TNVKD(F3(7X 
@Q<>?C1W D^6$=E'0MWI+NUB:7VD99M"A]DMA-_#I#&4 
@$760Q;<.(#<^GZ4X]\N&PK4W3K"^HPWY6_MJ!?4Y>@D 
@+;6EG,1+?=HZI[EUBQ<JEK%KU$.PAJY7OX,2.?EUWS  
@&(I(MAM._UB\,1X)1==R#D#_N#5U&8ZJ]YLKEJVY4.0 
@HQCBD&GGOXF"ZRZ;LA+](\M;0[X8IBP4_V%?QGO3P,$ 
@87%VM@,#XKDTAEIWU86(GLFT2Z$AX"M]BV5;[[#K>\8 
@&T5ZJU1@R$_O.40T 4!:0]D8=,T':E:*])[H(G+L,R8 
@J? ')32J=GAF*0\B!1J_OV B;'Z4D.R37T;0<$TC0-\ 
@EB?^<F-AT8^F9" 74U4[IO)J;(32\*CBMH$ULSUB=D8 
@'M$CQ>B%W8';6-ZZ?RB.HLWW(3H?4.TLNO9DBAF5/:0 
@BJ:0+9P&K\3?#(_.O?.O,TF#360+T4=?"MEO^;+%]=8 
@1?:T4TN1FT!S)-W1-_Y3=I9[<.>9)R1QH!4PNNN_>A< 
@E35,A/^F_+2426SC@E 9GHR+(/AE&,24-=,]SKW&9YH 
@D?\4QC$%YD9[L;7@8KEY+A:.<,B7HC:'OJ&Z+EDU1/0 
@3#3#:Y^W5R.Q[F;O'(VU\&*$1#1^W;T(GC/1VN:""<0 
@XAMID[&.QC4P>P@,O#Y-7R ]OP0E*675$,%"C;(DKXD 
@"MM#@BKO&,8U1<XW6;9]T^]?%#Z0D47=T4XC&1LMV , 
@- P([%+J;9_28LK6+^]8PM(NA0RCPIY'-S2*!Y;=$P@ 
@]:HR)U<OP);ITEK[96I0*6IMV,;6UBPYU^B?"ADMS\$ 
@Z6ITBQGZSP_BU8J!6[7TZ5 ;54DQ_]LFBU$3WUKFS4( 
@5BV*@%N5YD"67YGH5IW_J*(=,_3 4>R=Q[R2@'4E^:D 
@CURY3!-EWS<6@BA$J9LIUL/*7" :2I%2J:<4_^?G7HD 
@@L?$KIK)>*I(F.!@A;,A>"5T[R2G XIP]%VW$M8>'^@ 
@^2C]H^)3>:?R)TSO^3J.B#A HRT'$3+0@T/%'%*^LZ8 
@F,IW7<ML<EO-<(^#,4=5="SJ<>.8%).H(/J0*^,G?_0 
@2_?\81#^B.NG0GCHA^^;45SPGE !HQ?2[U*(QB-_8K8 
@0$=/\XGIM\A3V7[DA#A3!C8 L-&,AV8WV:#.2,C$5RT 
@X4%1D_".&1Q,<VVU#V!>@6Y_.)IR4^3J.#X)YSA@S4  
@L<!_0K01"@)0%R5&#)1U]:N304!#>O5)1FO -LA %&, 
@I?F*"MI0#/-#O^6G)P[&4+OC0>!%W/+\/F$?R0"?$N0 
@0$+3,#""P'&;F4  /3OP4._\P4C7L?&G'A&N!K]**)D 
@,GC]:-%P6C;O:1[DII 4%BVK'J+,/>A:& WJJ6@4.!D 
@7'NA50$16:UJF2]Y//M)AS6UJS@WFLA*RPMAAPS=I'P 
@Q@M>:I5\TATP%D_/:4,SR=TJL=&KB-%&DA ]S$-+HDP 
@X^5P-(?&?L4+PI?\)JRD)'BGT>F*)7B: XPNM 3?Z?( 
@'KB=-5I"7\:]"4L1Z(?_4W9\UJ PBZT+O&RY7O!$@9T 
@VD_&"GS;JA& %7Z!F<!30DG+\=KT^7V_*R.@&Y25FY$ 
@*WUJ3"3/KV!145H$U7' L?<(3C\VNBRY9"K'\(NIR'D 
@R^L"].W!6J'HL55D<B[K?MHWB*;K;/Z++:5NIG%7"Q@ 
@V2FUX,B<(C.G@^D$'?/G;^C&J@;_/PK*CE3$T]5E0LD 
@RF?D2"U-7=(]3?=3998OMEH_\=;'!-?=N<YL[PEC,/4 
@@15I#!EJ=4;35+EA=HHM0O&R.Q2PS&=>UD.^\7(])1  
@ N2$R482BRT=Y,K'_C]RM**QMK4;P-$/"!6OX5#=/B4 
@9U,.UR$%996%&>?>R4&04SK&:\#]ND/ <Q]I.<E8$U< 
@G3<.>ZK:8G9A,*,^96X!_?LN*SF#>J843&HW5\2QS&4 
@[<752I!#/T?#SWX@E,8@&KJ54CBA@DIZDY$'+V>TG < 
@A6*[8:,5DNORE;N6)@L8I_:@=QO38ZEEQZZ.[_"5CWP 
@*X 2H3M?TLCD__4\RRCV53Z%?ZSV_UITV1% H5J6W4@ 
@HHG &'P.&)_;!+!^7XH4M\V=_GJ)N#:XN+S#*"E*=,$ 
@GYB'C@MDMG6RAJH 7*(A<A.XO>)+)<5(J]KRYO'MQK( 
@2EOUVD2,U@SE^SPM@9.? 6T^WC#A>^41LZVW+9P!" 8 
@KJWU)YE@C=V KPS#W-_--C!V(O,'L(#=+'% Y@"^U[8 
@=/J\6C:YT:S06N9%^H;09_SACBDYEQI:U6N04[&/4PX 
@_Y6UZL1"1?5-/T_NA,"CCE#A[45..7<Y04? U:(PVJL 
@L;MK4.3E$3QVIEQB7L6I>X[3DU<7K1B+'^1!_=E=QQ( 
@Q]4JU--<K9HVW+,)<[QJ)8 \@<DP=;KA5(OB:_]C K, 
@^1/E$R[:3/#K3:/FQ10)K]R'&QNL8Z8G$BMFH8C/M,\ 
@88+A9(.<SGA5[>L0\:2MTXG4?Q;O<6(-R?,."S1FQ$< 
@W%O9V;DI$8T.D?!GP1*S3ND_LQ2UA<F#(173P?BJ<@( 
@L6L7WFP@S]69YLU0QVL)TI!DHO2Y*HW5PU<]ZBIPI/D 
@\0:VRI>M'2@B?D0R2S'X"?@'+ AO]I@S'2:IP@L> NH 
@T*X,(9QD!VM1N-SI8QY'F?@D@V/*DXU^\S*?+\.P0D( 
@_8RY,<+SS3F"/!N\^,V^N-XEG"]5?*<K!'F0HRG(A)@ 
@--#;:/AN:,XIZN$:3N4+IZKB6ZMO=$(Q<VNDM_ XO28 
@WCD5<OM4%8Q"! J<+Q:FT2L,]Q&4*']60"GK+' E=O( 
@;TUVFO.ZU%0XU1)SF(YJX/:T=AL.RKE.*$AW-L*/:D0 
@%8+H<^@H%4;7:.A2/D3E]43F;G^:8Z$PWI(X?1:].&8 
@"OYN+5D^YT/:XM+MR\6=]L!"1[?2L=PP>K>C ->HD?< 
@*Q5G:W"%M7#=>H&N6K4,SL+6'.S :$-UP2=9'#W-C4@ 
@;!XGKV'+-;^X>P<$MQFZFU/9IY&[C!!8_R\Y^ES]9<@ 
@*$B?FLC(UINE[PL">MXPT,WU(MXO%K^',ID^1]K2+RX 
@R&IN&EV7E:@/))QY^B"E.W,V56LR3;G;3-#3, @DW(\ 
@DOM#LEH?4J[6ZY3(EQT88C9]?"J+E&5M[$CV8A_EG<< 
@7?.7W_!HBUV0(LY>+X"3!%K[$KPWJK F^+612AHO_5$ 
@83AK@CE(CCY/E;J7Q4Z5">'3=K7.UK!U!9%D(Y"#<@L 
@2D@@]296(P>1D,V<,#!L,ZG%6R"<()&Z'V_C["Q=5)0 
@HR70BIOB-_ST>A V@7GKW@")MJO5O"4D0YL+E<:REG, 
@%H':TLCNPK7#<\,#:O%AR"'O21]N&6Y51.GL6W3:]IT 
@[@Z3E]TDR[9+HX@Y^!N4KC]QWN0<-10K#8$@MET;NG< 
@S@!6G--V5;CN\"67P=+RAJZF!;!NB4AHTD\^!BO/ ND 
0S*DPGY)U3HE(XY8'U<&),P  
0>452OJRA7D6^XVO9K54.HP  
`pragma protect end_protected
