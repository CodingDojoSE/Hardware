// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
eDQDkmfl9RuBPN19lpm05rfmhsJFIE5vlEFf1yWY1SnLYf80HGTL5PkISWNG7ZX2
d/TbuTvi+8Q3WDezOBx3Lkgebm1FceoQSRX80+vsVrWvJd5ctwNBW6BiF0NjELkR
Zk9mLCK+EQ+e2Lln62ilK+0CE5BjkwgQJylCuYD33VJt0kPPRqod7w==
//pragma protect end_key_block
//pragma protect digest_block
35ZmiENo1/gsZgUEUtrVHtkiJQs=
//pragma protect end_digest_block
//pragma protect data_block
rJoizBBogWY0MKfFoDaqdy8EbDsU7hfhZNcb8r6xXqIpheNR/B6d3S1bCxJXolFF
Qv8gC254JlhHMaF4XWbckk8dUkTBW7O/2JJQyebpTWxESJLIlNHQffOemIZN4S7L
3XQCVZoRrME20bmJ6VyiRAoVFtVmxA7KAA0zEI+4lGtZg6X3JG6wGguWiejnakXX
Rqoh6aLKOXbneILRPyDyJzhiDfkOs3m6nbGKipUb3bxKuTLGhjoHuprLRpUDgRRG
4VWB8qEYpbttZ4AB7QQk4HHz5tZPayq4iwjkVf50DiRf1VtaJep50SYMbQeNCJII
4xGlCCqwMiWq6Tym/hfIk49d01VKJk6pJrEgJ005gl7X1u8o+/Gn5CgZRqn5bXqO
RD6/WEgOTdOUaGqeQKyyEdsVgwDq6/YVjp+eFC5dxqxXZU/XvmBctUnf9iwpnd69
y9BifaVubddIFUHYKvOt8iqcoQ13yefR+zvGsX9TJkoUnJVUDxexMsUeMbAvb1QJ
6UivNkBiNhptiVF2F/l8kC3k3mhurY6y5w16ujI6yua1wUXKFSjARPCoIKh/qhm7
HpxMcq+WzETryxMWTvuyfrTK4wZf26qxjVY+6mUim6ZCBUTNVQhWG8Mc+SA69GHM
I0FO6teoXwPujM6m+sklzYU72iM26AUcebAWGDClHxgfpf2vVE4m38q70+RHlP00
gz4QXWb8UCJ5OK8kAGYL2fUxuliw3G7caDeBDQCa6VjClMS/dLkjdIGQPb/ce6eD
CJKZpbOyBI3FkcIAht4vGwrgGixlrH2Q3/Kzya5outNnoQo8KDgU1XnKGvv3Rsu8
GZ33Y+/qej8yyXapJ5synBw69bdLXxGcoAbV8tY24UUhktviEi/1NCxvG/CK3YcF
c1HAwYbNGk2dkHaID2tD4BGxUb5U4mAUL2O/ZsOkdmn+IwV0oENgipicupRJPC/r
nnxqwrYu+1RUL//NvQGlXkb20TjeoCPRl2hEP4148bFa4J2zlxrjN8g4CLhWxYfm
BOEpzaSDU0ngILAk4CJrmZYjV3mV2gp6s8JOA+VsInhGHcQ9Cf7DMKpncXtsmwYL
KxoLin1T6VZAUjyYupdIgJ5LwuyGEBHvVnYYfURNr96ntEMqEVcfAjB3Cu0kXEzQ
xnyQDYsLI0BL18cv51CCaooMQT7C5eoDQxzJrCTk3ZeAbcCZ00FI3ti5U3JSv9hh
aVmSZqu9VUPfJhBx3konuaTQjc4OdFMp9Su5fiwSa3ngTuA4NDATqH7Adtnoo24W
hV+qP01ygwYyGYOyVnfcLphuAP5Egeq6RbUSP3OSf4r7lNghSKGP6AFXsYY8ki7M
jkYfFlG+IvXn3fl4DliwW3EwDiP9fJzNH3iztkX0jKyautS/2yI8Pkg4gXyCCyZf
hxezcQQG2J3IEG2dqia5XEpfr7cnBvGa4UYvGMaYDTgrNqNsChffw7W+UaVXdVq9
EdvATC51ZnOGU2M81990wtANPz8RarN2ZXkkkug1koUPqGoHMceHUIwZwau5F4Bm
IxCk5+72Y6JdyJaSb3esVRNfuPzX+0YgcbiVfHwBxmU384bacS40cy3GUeCR7L/s
cq+YTS/nJIZIpiOVVk7NpOE3cPihYmy1Quf6aOC5ZuRg6x/z7G+kBtgxiyujrtSQ
CqHFGbEU94BghRamGMMWvkzUmVRwRFyqmUzS6K8UqEiuZgTkVheBAEQ863DLomXA
yVptkeBRbfY2WzUaWZgC+Rl1TDJeSx7a3j3pJwSjwXHGFFcSxlJHlCXj7RWYW2YM
pnXwOBsKokD04jOrWZyUR+mC4bMXU97mLYpwPM6vL22C2OCg2NXQ+dT6gTiebxiF
QHOerDSCnyWOZbU6wKOTk9O5K5TmRoEO0qwzkdp/FK/h/wy3n6dTm3DiQ2HX7uDn
2R6uC5JXOuKSIYbcygVxg54kKHsqjF+2J9xpoUmYBhnVHi56RN5H+9uYaNd2qQZd
7m5Y1wuWVrNY385LiRs/f0Ir6FH/THEHydZOSRJSfD/9KLKqzHoYB8v6sBfHwkxW
M/+8xUuR1CzcUIJhrnQ7YcURG98Ty5EVXFQhfsCCMYPgYrA3W07eq6NbIuaNTjL2
uO+4nmTlkMdO4C4p0NZRbBFdixEKPhQUDBs/RcILQHGbG8uG1my6Z5EHuJre95Xk
M+q3NG9o9iBcomzYPUGjU8dsQuwyvLENsgmymYIHMw40pZxKDQ5TNA4umYsZr6st
FcO0Zh90HpZyV6iXPIdyremXkBHfqGjQxXioOnN04zMnkOHIZbkaBt1sQAYfhDUu
2o3kZJAYcxPW7UDRdKyml+kwGeLbYrAitBgNUH/sULTiiU0fLyTTs9Gn9+6TZwNm
WkhMMTesc8dNx9KDytF3394NVgPjAcIGFYPdiAdXdFxXxLW/YhIwjFM9DnPRYMEO
nNSZeQFKBORwsqqffZTO2jdgAwrWwOpLZ/SjVkEQn9Ia7M+Xz0rfUDMDmnLOFFLA
ZE8il+VEe9J/y7ZUFRCgkaCq3cstr8hQN50jwqZOeANGHluhw2OHgYOWGoqrVGmp
ntIZydT+vc/9Ig4ETwutpt+NhthHvG10V/uMfr/0mtH5P6RVRD6L5ZyigH+3NlNR
LQMofqoY4vW2IWvOESXeVl36DXQRbC3RbzL/XT6STxQIViW8ocaJTN8/hKhEWKHH
xHUmFudY4GyzytLmDbFyTu13VMgmbAkpczRfr+Kf72qa4hyiHtNChgBJVMNTvfrm
XPjDdpbrnlkv+zu4PGKR12lDo2XwfvlWBZK+QQXKABlZByXdJlmB/3exwYqpl/uJ
DgTegSnMdKvUKEne7kj5eOjq3t9Ir/oi1m4FsoGWnt/he/nFzXLLky9eqaDPxzY1
Jcpt2f+lgVNr+dAaHEUZQg/XH+dwwaULh1ZJkTn5n7Ya8gDi4nUV7AXCknEHJF8m
zsLOZ0ekJOvrKXIrsrypXgyvjERxdSr8XkdLIHERlataqGHlFZCzop7kQ2jgr8Q4
9CokrseqkS7DQ/w8PAl5PYg8Wz3njgLnlXzrQkRxaFmcPlEg7FLbqQUWTV1hNI2O
dlFN+RhhLT69fDLrXlJs/CzBe/1qh1qUpgSOcnVXdfJQsMOU7P+lpCSjdQGOJy8C
RJ5MJoKI0EcFtM4zhXm/cuwq5GC1zlkwcHYkSb0VlGgnY6ot6zvE+JVajDh4Y4Of
hJY7lC99tx8EM9D+C1QE1nKNX+m7BExTHSFyJXHHq0iBp9IPnpYbE3TmjDGwra83
8iSuhfeeQBbbAKtZojf8s7IaR4UYAo8QuFgfdU8+I8nWZftiVcdJQ0KtTg05Ff1J
4PUP4RLjN31amxEGBypGNGmF+DdIvujlmSn2mICERJfB0quEJivJpM3YgsPIUgvN
1xhjQ5w51QXg3ZJPtWW2KsLf7EfdWeZKwEQ7i9ftBQV6gWLDcd4mP99XLRpmLxXz
1xqQu383oggkwBe9S/9NShq+R7Lm2MAGX0K3oGXPpobJJ8CJSwr0CA0GKsEo7K8q
AuqixZIPtLVtxHb86gZUJnqc0348TUK302manVUVxxPgGvuSZnD3XMl0sWUNCW4X
uto5YRsG5lPQe6XUn9iHtkbsqhw36e0nVUKEwlANiceah2wujasuOqrZJr/W/SoG
R5hWN32lxknJTrcTtmrpFh4B9e/zu2uiyKMUHmbN/SAv9RwZgpfwtzU2cnnm0q4h
kzTISzy+7aGX5A0OBU0G3IuICH/oOqfnMMOC+LjdX/eLagKaVhipz3y3pg3hW88/
BCAFbI7JfOl+1/3xqUvEaGx0rVg8fSuRFjFBzNTGG1UYDwCZ4IyyJq2X6hSjBoES
Ds02Gy91SSuRH35jSu9Utaiw0l7m+p0mfO7CH2Kb+XdcLu54rKb4t/dBCUw3QArw
vu5k3ILKyZOJbkK95f/UizmBjcEODHBtkHLUCkZpNcb8rNjZqQ+VYNbLVzfiPheT
7hkhvkZ0lmzYP+UpqXQn2Tz/vRJQjzL77h+tNQZqD/Y/flIDC626Zxjmcp8R9WO1
PA1pPLNdw2/fuWMYsyM7BXnfL+0S+4ZeIED8IUxDOukuPXyLD+XZz4MYsNWx7JGu
YZNsbQEM1CaMCHgVHljR9QNloTls5kXhsXloy3LUO4nZ27d70KUCQ4HaLp79EGJm
Z3xtVZRaguLdtavO696n5I9oMgvV7+TbOBOYt+B3w4cEQNtSgQcumY/TFcBvnQ0o
L9RxYNbltciUcSjbRdWTp4+GDlvmsmL7hf2tGTHs5KYwNa93FmzSga3tjYqU6gha
EGeQZr4jsT6zIZJFzDnY3DRsb9Y90y9cUgoTNVItPp9c0Xh2Uy/X0/X66pIHbTKK
j8gcgfLlTdcJXKbV0Ba8HP6Rl+nwh1jneXkcFYnZ9LQwPdN/B/y4qkjd7qNj6GhW
4fbW868J4ez6uYXfin07TAMnMhYTD5kohuOWn2QADOW8WO82fZMRdc191UOT+Pbg
Jy+hbQ7ATGJ2SPfyFieukzgzJPb2jBymg++BISZMX+iQxA1vWAuVbAnyilrpuu68
jw9A3I32jF2dn46AzesFp/cc8t3+XKG7vD3f8H5Y5RtYSzGvtgS9hn/8VRB/8sbY
HstBpI7BAHF6216Bug23VulGUXufe4am5vZGQNtRCs/dlfZYOqnLAqXgbesjJqWU
z8a6B4NQY82vSY/R2epznC0ry/+HFOHvklrEXNlbufiM9YWKqg9ZnMv6rhNIVZOj
o2bsn5X03NbeqnOcVS6TyzKBavjGJYM75bom5px5MyarIao4eabdj6vnyYzn6y8P
Yb1Rq3EeVYPSoQZ3mXMlFCH5xwOhh9bMwdQtMe82ojX+1I66Ez0LA4g/XUIC4The
kjrN0nltsyDO/nLKyrQKS2jfB8Qz7ECXH2fkVRJUsA9jETTT7j9lmpIV9ibMzw2m
dudhTvIE/vplCobB6UZ2h/eHEbudZyVFQ4FVorGTZR95wcQ8v0yW6epAcaa9gHqS
hN7PM09/xN/H12uvcZzF0BgnG3LXJ+dC65MPCFBQonS70kG04JqslVD3am1UCg8j
LJ0qISnU28TAIo4P8wxY5OQ0XNneL5rRRQp/ioNsCQ0XpfyTjxFr34JiLONqRe9T
+7lfcEim/kmE1j2IWcZUWHgmpXq2QYeBd/qGebgSPrRrz+WlsKO0Ek4rHkticC8t
J602KG8DAon9vZhN3md34UZsjMmP/Nr4nb3m7cjZ0n6G0wTI+c/yU15Fleq0QQBu
ZICgQgV6uiYJawkUkKgrMqA2MtHC1dzGJuhxskayJbykC0kOnIicQJhi5NTb9NWm
Tffb67ntbp+PefddRIKDisTfiTGWAZNCX8GxFhznU8IvLrqG4ab1xECMzx4XjRtL
Ev/xwc5Syhdce94wbh5hxAUaV27g8uo2OJ2aCQ+TRUghBGhOPadlKRBiSZvjJzY5
T/QPbKEJeXiYjPBwtSQlYqDlNOV+PsFdzXYNk456cllNmomuMqOmOy1i2VLiqsxU
3b7slvQ28fYdNOoWjJoAuZ1h7NoJR12Zf5A/9frD+Kj8mZp1uAyJKsdR0sVhjMc1
Evw0Ldu8nQ2gLRTTMBaaDHA6TBbIdVFVyxs9GjhF0bTD50Hp8W3wHIb8i6SqOJFN
TMZK7DbNvkpv2jHGHP5HZ4a7bDrEEUnMuOeydpEI31JGyaHfMAic7N0x83XWZOT7
wooEPaEZlxGC8B1uGhYdBTXs8INNAgchjbMpyKpiRvJhgnkEwA8HnEh+FaGioay2
MqF/lH2Evwn2Z6UhrezUrv7h/LWAEaGxN5xegORb0CuHfO5LfqZx52+Jej2PhTOZ
1ORc5lNclcPpQJcrf+6gtZqpV3L8zRuXKXEhkNjvLpYIrMXY/CWgn193yyZ9aXZ3
fiXa9/vGqF3gp+9T9cL08yTLbCFJ6Ny47bQvCPa7ri2QBLhZBL3it8SmcDmQyZko
bc2Miq/H9FqmCAffiICiFVkRd774r3aIuu9Xe6mTqAyg9lWiByoyBnAiLxf1yXKp
1s1YuNZhUyLbWlpHXsKxOr2GVhH/01R7qVwSUzVcdWw9QHSd6i5aw34SmuesMTLs
Gi9r3UbXk8dhEey7mjHQ+hCJG7BLj/WVanCmaLctK6MxVCb+zKpS4dabZDIkpqlm
XIEfo9hcmcemQZIGnTzwdPFeyhN22nx5bVv/HOSOkhVfIPCBXhFQeD4t6TnYwMKH
qFTHVw1Vv7HbSHzzpgm/xTqQBuY/LSVw/iV2bcXGKKxvJJ86ceAive83imegRnP2
cYDceyELtPjF5oyqYzpyf5y4RzQszGv7papGIJPC6jDrFUXNq5SNVSC8Sv4JUuvj
RhzlpIVWmqR3mrWR1BdhiX3xpiEVAvgbXVMox0WRj2banvJ5L2NOQliUqhWSjva6
zqe7B0Hgp8TF5M86LS5KtfxQ01wAeEGB0MMgnhxghdiAx/UUaXd4Y2al4OWjHKu1
2f+fFPB4DQ8z8Ka2rzcrsEPRGdC/POTtdKUwun+A4mR6MDYlCj1ckxKhFO8sQk7S
7nbUHTtj3NY10xEDbfM7nhOPvI269Avvu69KCexyulnFjPUBnT8WEr2vTJrq3c02
UHZ1xYxH5Q0I6IV+6pG6LetKvk36yx6T62uyRQ/YCmtcrmzzOFhdEmuhHZHufnJC
7zOyAOb+es6b5G5JU7cC09CbDMU1WWxKodzOTyyQJdhCZGTCL5xs0jGU3TYU7xmL
tJSXkBKnu5KcmfrncuOtWd4zpNVWpGu5Wc0Ti8kNwfEXJ5Te3MMwhrWXR2p3gNWA
Mmp+anuAOclI942V7YfmF+apjED0lOP1fRdNkE1ZuIOAJM3ELJ3AApb+fqqcdvNX
QFf5Q1vujzdHTDLl96kQNXQ0Zq7TUbo/ne4KvAZ2bY7JdsxrTM2lQ9QDY4yE9IXK
eUrxc5JkXnknv3i5PMxLIUwEtx8NgdxDC3CvExBTpA7zLY+f0hzZ6bYvgMMuFZ4u
E5QZyegs2UnOx8Tun3lHGQgt7httpqQBecx3k2VUBZvdKqiLyj+etynfiL4l4a2k
7w83yBuCH9YBIVMDAfvmuoij72NEaZpCiB52pdGqVIumiNzUjORuz2T2i7XwYHUG
2iTJh64mgFxIJKFF/Is1w/PFzxRuLEFG2b3GjSlj1/V5VtaaYc98+wHTz/ZKq/2+
F55t23vUJjxX9Lq7Fx0PcyRnfwb7FeICp4C8qy0dUFs+DOU5vDDk+vBKG3Ke/91Y
iuumqbu2dMLAt/m+sXqJl/ZcgyZpfcQi5hRYpn+t6cjdl/0ExZLrU32ZIzhm0gJZ
RAQi/ZMEiac6wXN5lqXjl5ZBOQJ8xokxnBnYtq9DEgiCNkurk2cdeoPlmpPzDazp
38T9cbMXVElF5bXj46fxSH3vvExhPKz2bhlDsmP15EV/kei+Vd/pAvlYSkDuL4+D
57azS6TkNjQ7yy1Z30uWJB2McDuC7y6A7+WlJHcQlZNKe+8Ox0bf+ubhnHRzxQT0
l+ZDjjf4EfgekBV5KsVJkd3aqc2StvWN7RgESVL/UNKIWdFzjPpHj5AHZ1tVxeYF
O7vvXultx2iuaDWpGG9giPyAajs/TX35FAAvdzUU0y30F8U8vH/ryTmBsxiQ53jx
nPFKSBVaNvbasdH9pcfHLueddI/NmO39GujcVb8dAjMdwgj1kXyMghPSy8YTHc6P
FCCG6AGHPtbWCl5gSDVQ9zsj0HVQwsqmKx3mFPLa7VBCeCLgz+YgZoZxnhHO2HdK
3tx9e8d+/ANphN4alePDCXb+67L5FwGHzfZT9gg+EtmPSC4MprPVQ27vj1cNbFRs
OxBYZtA4Y8F3XSe9hK4ToXDSsWSIGGyH7C252CqZlqzJTRo7nebZDNAuvQ51sN6P
5GruIk233hNAccjikgKeb2rRR6c3JooMnBIVfa8z3pEuXMR5+MLYn9Hi0tvNVSFH
gNGI5HiuVKkqDBQ6XqqPdAPAzS6/QgxA9UILaZWs6bBEHKaUwcsuIJMQwsYwBHAv
+zhTfAsgVEUjCVbZlZwut5ng7ozHGQ9MR1+H65jNWRHQeVdurVSGsME7ukiSdTpN
FLRwD/ZFIPRfjH+yVeOY2lQdMH2nL1CiqpvXOZcnBR9INTibHrbKkUVWD6lmAoLZ
N8Ha+XJ1dm9hBmdLwF9/gtIa0PgJDxM4gZOaZ8JDHvqBIFY9ZyNYLizMQWgP4q/v
+XVJO8El+KXsY5N7a3nyvq+DjnuhHlTozkszDYnKDVKLWXpgHZz/nwJ0B64pqHv2
mKnABMFpd0eKfndyxMs7z6lczSSzuIfdrobVCFOlMJMwTL9uILSce3aShIs7d7L4
AZ09OSFOOQPC3EATLRje/7WUIq/AFSxbw6o2qO4esVAlGt7ppS5ILMpSboEeNnNU
e+z68OzsEv6Ukjl/TlsaFZ2dA+/jUA7MTQeOYaxHhdzG8v/BaoGZuSDsUdZD+yPL
Tsd2yuR9D0Oi/5OndZht69i9ZmB1jsAJktjmkQ5ZLACawbymNiUJ87N8cyDV3epl
z/a8juVdwa2oi8XKQtUYNbZYZDUSAUC4+0fY3AogAp+HWJ1UwURKDVOOPcl2/PW3
4Bjh5GvMu8Rd6DnTscaKHCTK9T8vOZUzp8L0vavcrGxnPEZD+H6xjL3fKcz5u6oZ
imiE+tmbANUE6BYBU47moCK+fzS/ptVOcsMvpOErRE4u8PsoBW07eFxuny12V62W
KHG2SjRGQevxKuQMi9+RszlEEW1xh/19dVrSVZMQ1Ndzug/WwupCnzAhoehYqBBw
FwOQtABFPaatXL61jce7nQXseRPDdbg3Bj+aKzNG2IDmUVKJbLcNq9fyqr9oiLvH
Wf4wsmMkpHzX1YjWAKx/PHcZiBlSvYODHjCsLrV041n7FGCPZ3w6zHhlDx/VQVdp
vHAWrqRKV42DqbvEmSxhmKGDaBua7zEoxxVS0jUdR/JCGUJyUiCV0QngJKyg55bo
/q7E3orRa65LJ0t/u4QDb3kF55ad3qs+Tc0yozRGM+3pJHlta+i0d2lL2uks7VWW
dEppscmUqdXoePFKN0NkRAE2ijPZvDYod5Q6ac/h7KXVdWhBXQDlnL1tpy3ugW9B
yOPimXAC6eqePvpuq2GHJ95Il0NKLOA7czN/M4e5lvL+gNnMTuNj9WCbdfDWXQqG
vj+UhufDMH8J7iS7rNTIhVSZYtBWum7tNmStOFRGCvCNhOVc0Tm6t3N88pF3lAZ4
vVGIgRLthOih9e+qGwtoJAT7MtqmzjoBk4QVTRXvqP/Sj9bl7FmnZO8D4KouZIHB
6sqQtD0Pcl/pAHX+b/YFR6RlVqPfIxDK0hn5tadg+yu/lm4x8HeBPY/iulxoeqNQ
u0NeOsIp4WpMTAgn8+n0cPgf7Qe+DeqSsNlStZBTeSgTEi4FuEdUWGeffzCdIzGR
ni/2Ap8+4u6gde7H4RrOPyE327C7Hfd6K1dag9tCXlqU2vvaYkO5jZGiyLE3RDDn
K3eLDkBjxiShcGJXSJPTup60yv1PHHwv96ND9g83jM4Shjhq39IUGexFDqWVuVV/
Yubzz32fHD/0QswS4hbxj2G4h/7C9nY4JmS+CR32f30zDDxp94KbHCUstk/GOQM9
pyPjIPR/1HfVjsf+DEmxdZvd7JnNKlulcbRvpJXWyeqZFH0lWiv/pkRNZK2cd2St
+GOU9u76v7tKsKrvhLgACGIAjSOopUez9N9pnI4ZSchekMOGq7YxbSI0nA76f7fA
NcnCNC66Z2ZkoJpRsT2wyQDWFQiVH6rmb1t8oHgX+wzB39pfWle0ty4V3QVIN/XD
BXYXUAMju41aDjtVYHm0TLQLwiG4wl7nkRli/noLfzL7ycUZLRmrK7s7ntTskVSZ
ZOPh9NPE7GSSWsg2o/67S70GSstCj4iQnePhBPZz41RJGFaxAAOUvmXgZGRuQxDn
5bGlpCbpulT+dwmtOEx9OYnhp+FOncjMLscYZ5Q7Ci1kb9HQuKl/JytXSWNe7tIK
jWUKaxKLTC9R0Q4aHprPdqAIIZ20YMmXhxHDgP7yZn5+Ei35xrwim0Nu/Afgj4ps
N3IZusH6w7JzXlfCIOaPfvX8EAThL7gYCNhIXBJHes/FEg+mS7SU6VOVZtOcRQfY
7br2MRGpm9qSd8t/1rdBMD5o+2TDzoQ6+VSCuSjv1JqPC79uXGdgVLeCtfcNkOsl
Jkz+jIFRXVtCbqiO0/g+Wvzt0iabxciij19ab85NrmppHp4yBd2FK6jiSPovvy83
5BOQAmHbqbO8SAXTmX8U9vgmbi870IThIIwwl41JjqJb3rUCdaf39VxUObhDAhqi
4/f6jvwqxOjP21AF5c6s7/X9AqpXHGiDstBowoHw5FEos0Sd4hdPTHzriZ7srnF2
Qd1wF1K85JL9XvHZSq/ZN0BFDHdsbvfNXuNIubI//PwRc38dmMbF6SGzUFaa2LmX
f9LSrOnXREZfRE4qjlrtBQSJOKARdtafquoxofT882WuWGe0zDCZgUDeOFkiDPDi
+kUZRKfikHHDoS/h9dXDeciI4TsfRCriqjoHVUS6rZI92ZijbHEPbMQVTafLHsG1
ORNt/6zqPSS9y69KLvdfB81xqJQ3Fluh36r6Gm3NH1beQD9XVNlGERlmKVltWjT5
T0KhzYe2/wjAT4gYzGxnq9gNMXib4QOp8LhYzEY2npC0YmEHyXFg7Nc9PWUfZyVG
MotEcAR4lSUYuXIjzQqgB+W0MSluD/OL8vR1FBYjLjvkhA7KPH+x9UZii1eSxiXJ
6xhY0hYbWwdD8iecloLqxnzLfJl4iwSPJPdHlxWczhkEt8Un+UpAuWxA2gPikL1Q
tqylHYCfu17YEgDD3q2jcd781Nrtil3ulM+2oT4iHGiO2RJS81V/sl1Uq/u2NipQ
R7E65xE8qvLPbC1O1CwRlJnjY5tpJAnjCfgIb1T38nmC5bUxVr+lNa8jSeuMJyT9
29BN9xTVQxrvOnJUwVQj6KJnkl1VYGoovOriNONx+hvjgrFq6hbTADgOTAfnxL2p
/O1Sx7ICb2Yzof6Av538nU3kqFYmj0XNABMC19TQXibBiL+NhP+VFecKx5gy60IS
qfuyOyrujCzOtoITESQvxtlcPmZxKDlGTLxXRKaccdcjjlqUQjsIZcp26Yx5hnTx
lLfFT9/6+XO/Ae75vpOyVh0Gwm78FS04SH+09mzdrhg7Fa9IsvwuNbN4UaUvbVtH
5kgyiTzbdKUMfct+LGmij8A7rQFczphoAsfwL7dH4box/0QyERFDZutR7GpHV9GR
CgYuw3TA6uhe2LwRBVMgoJPATsXo2h5xTzCIgyPkHcEf7oDcTtnOgZAp/yq/3jdq
FPJBzgzhfUZBpNNFVZ6xMngDnLhAUnLIiExorkEyCLweyADlvh22JPGOHNNmh7cT
mI/tYlnKclOSjEmfz2cYBrcmMZ1KQdloGg10xtBKqgiXmmLos2P4RLANPL3RwxtQ
GvCGD1mWDYTLIfqes9E8ajA6sFmlwizHXOUj3+vP7xZujVjyB+iIWArgZrv8sCKa
VzBm4tWUPituLBdMbx/0SQGjswjz4eZxhVRd05ZNT+vsPkH8SlAiWYgWgekTzYiv
c6ZixSvfwzYlh/UdvglCdqYMFG1m9RWFQKF+iQL+JPWX9cJ/t8DSWQ37INbOuiZ9
z/itO09XiJIyIhNrWUed4Jl/m+rWzhbg2wq2HFev27bOaUcdr0eibHPYsKux85+2
RqMSn0WgEH+sIhLQ5js4NGjoFe8BYhFK5oOekWYS9xvKusKEep1NRpDa3e1yk+BN
iG5a5vUbCLdDd87mQF6HPqWqIyESAYr+9K89jblzOGiF5S/mb7KOnmkW+hduNldO
QgcHVX0jVjwDuNhl0fU1/py7/l69p9sFythvdDlUwkCIFMG90XXRdFFgDK5nqqMQ
9kJhSKL0zZT4qoQ5/EPA9Pw1OBef/M8HFrrByMIVaRkNiRWqAsG8qQunUmQdBhTi
cDUH4lNFCczlULjk+7/QzhubMBb3WtGaML5Z24K7u1nlU42ps7YyEeZUkPsu77Z1
LxJGYZG6if+JT88u83jDIXUXZ7NZYeKgJ8Ooe6XqOqJ6Mp+QEDmWKHN2ZRe2hk4y
b5aDh0yzdkpLhxb/tQz5Qaopzd77evTfZLlCabmBn+l0skwtzzaS1of6gSqte8Ci
ajoBH3HYI2R2Kee+aBmE7E4Xb9FI1XyPQT0qFqjNJN7MdsVSEIM7b0czV9ku53OU
b4cnVwbD3/lKu6OvnHjfgmGqPnCKlqqkofDTKVMbp40kZLr4eTa4iTUZEbTHQj9P
q8V+tWgn8njOntbbFt+EF/EvJARTtGVQMIt/6AUee7N6uQODIRsaYdrGQ/leD3AQ
B48kmMCoPPT/m2CYRAZwO6OjU8+1lMSEA495pL0pEkhhRFaX+gXgjf/yqnUZ6w6E
B9d0sSQ62++5EUAZ+l3oUDhOrHtNg7fEIEjXZbQxUSUq05TVMeL6Z/VjtAPfN+Ut
AHn/LPjw8Fsya9aT0Bmj8ZuvJxmHV7D8CZZujca//W+INQYisw8aLi8opcHfZqHu
NVKwmyw/+dmyrX16EGCbaThab/aahJEG9PMlXfBmyah0Pu523tMjlAw+bthLRrNS
wLs6hNVz0LyNOa6EDHRyx5qyNbbfFiuvla9IjEHsf1qxEigcB4/QAQu7iTrnTkjs
vfl2WnKpyUxTh92wS3wggneMeXfXk97kQIlCV2wvbIfph4gH0pnmbKkRAc9p5JY6
hbdx5WT89h6KpG5zLGScxGs6XfRRyTmb0DPMDYuxVWlu0AJfF7T4nniNNyNK+pMo
+vhjcUIQKQyGaFKzoS1XSXXEKfNGgz7LrKhZT02BViToZBw0A7a2i+HdHrBkYSNU
IO3IPC4FlzbJVJ8aRe3ZG7PYYGAR0/Xx1FSKzux1Som3n3nf1cFr76ZWAhYmtjFf
sH+cYSVOlFc9SqOOyziIMIxvEGJ9jgVhxD3U+Nm5daxwxjAnb10P9wJHVEb0cGWH
5h44ZcUt5ndXqDRbwaQdrPrgbD+DvV7A96E9PbtL34jd9/zPsquHHd9wu0bi1eGK
SkRUOirRZo9ym7VjzhHEr4+7ul3T0BOkkV2SHATuZ9ybSmNx+SeQUhQ0yBaz9mk0
cjBKl0MpCEkXzsG8KPvSJ1QgvDlIFjJUKRkhnMUpkoUFQefuC+lODyY4riRhBZtK
xTm6fkRdVP7gjdy88/g1y7ev9Cuc5V+Kknm872StnMOXd53epYS15UfLTMFPVSGc
raaiQMxH8WZlsq6D/LPmOi4+JSJXpB9AuAsZ9xthBcYwAS/5Ylq34FTXaG85vM5z
4WPF8pmlREVMbdvpv2iP4BcbPnuwfm2D+7mzuzd1ZT1GQtbxChYfiJ9cjBexqj+0
3MT5rb9pC9fy56CKjIXHzC5UUmS1muLmvvgLZyc48llTm4uJ4DZ89qIXduFoGOj1
ap9nkfZedG0ZAvPQd4c/9q/ZU384iJKNswt0TOD29+Iqot02zcNTLlkB7+7KcKzH
4+fUNPHwz9xx28gKta9zL3TYlUIb6ANOlBiJojAiNlgrxXyZMz4Wg8hQpBNfxeLs
59zH23MRiPk//Jggzmwr9qSAj2FRPnz9lPwklMwOgrBODrRA/wxWuy17QhGu6+zQ
GhX39e23q3ZgKEwd1yadbJORjHNUjdx5T8KSebCPSaQCCAbhUZz05hk2Go5Meoyq
YTh6zEHhao8rYhGjWYjxXi63no5gNYRYBO3tUQVuEIB4HW/o7qv0hdIsQqef+l0n
mQb5GhqbDWYbjqGYxSVNKlHa96omMQqMjOiTurJsWYz6TkjVrYAqkH8WZCYefBiv
R6xv5Ys87KcX10K5AgF4AWBTZBIAQEB2xTY7WKDKL4ffbGb+TpWPWnWwaHI5GuI0
ZisnSuVoGQL3NZhsBez5IKQqKozW8R7PvGX+bvbcly0337w1I3/22DdNQ6+mkqy0
MbTxgiViNtaIxgGXwxLlvxN7ZndmxlBaIv2Cgvmph+dHe7f/c1EPskFHXnex1ZDZ
xtA/OEH3Y022peu+4Z6qJRyry6BIquNvRu6kpCiHu0vhEzHXDhgHemG4f5ufl8f8
txVjkHN4BMb/Lzj08pMNsYYyXPaP+LpkualSk9kMC+0R8HXFOHLBVVVEfHEkkOYi
i8BcZ1usU3Xy7ac1h7+quqi4snluOizZe721QzcsGdPrrhHma/Cvy5x7y+YsHdDr
25uGEFoI/zgHaanpzsjf2jvcPSZKkeLUTRKTtcarJ3HMU/IuABO3DvH3ChAasIqD
DUUuwNQDFvVbgUi8Z+gfiwvvLuEhuq9QeCVt3NO7Oc5g5I0wydSLNzXWOCSlliuz
seNNHTPAEh+eZyW61Ldhx3/nz8wBB8euqGYWnZ6L/+7YWd7kAwlJqnzO40ihfKPT
NWjfIDLWSbaYUS1AxYLfX5n27q8fXIWzyZQIPqpNWdzO4DB+B7qDMiPLyYdi3BGk
itOM69w45wb19ieKXxb2Ux06tAA6KQaTMW4WvngwjsQLRA8OTwf/kiSvkfgbA6oU
jduWNhOtbA+e8QS3CiCpo+b1/gop+4KzwfzYBBRNlUrCb7jZ9gIXtN2o5BUDnhFR
+JMOkSRNd4lco7PEE4kvENM1H8ERUpMtafWkHYHjVWxKqkyGFGqQP7MFJuK0zt7L
0sv18vccI6/T0asLw78dkPvXrSfMOHDCrMgv422nhLvF/HNexVva3fTH5X5bKBm1
qG4Uy2mAO+EE+RtJhfOIyOWEneB/2w65G9ThPiSl96uJKOGs1ivESFuDKRyoDg2K
DonzF6IMHdn29g8tqcoKluSq547Ux1BmbxNRPlMPhGrvwjxuN29aRx4nILArf4OH
gMP3wuf4BUHHWEUAK3eUqqQ6gBH6TfLJ6bUr78Ak+4ooL6AGcblA4jbvwSxr2yPo
NChCAMjKw9+BF98Kgj4dTngiPnva+mVKndyHUmzaSIc57RE+VBZbIX4cvEVznd9Q
PJ4oK/AW3d5p8T5KB5sY7c8R1wGqZNe2HgoBLSXbI0MCnihlbVdeRgxxnNljCXJ6
aYDElw9f4ZI5fje7wO8+Mzy6/lKezqXWOk1PpZwo9852k6Ve7V27xeUG/zx9P6VC
O1OG8/MnE7UTdQzjlgNgRvm07FmfGJc/EpCs2s/CcDimBLUmIfDgZ9CmptJq+c+h
R857o790tLjyT+IgX0ZYddzT0pb7buDtSpONFnZTLO6e8OBWOWUXBSNZN0lzKovt
O1XMMn7DBSvf/BNEiOpJe82GC6ZlZTr/7ymokmUq4tk5BncvR4jXw4R29ugENWRT
M2s9YSV5b1KgpV6iIpdLrbDVAYHwuIEluXCV/DaqVt8JLZqFGnhapPIt8v2RTF/y
4ocFKZZ38xbLlCNbVAsrwEmFmpJ7xuuAHcW1KFW03e/Jyc0eSemkuIRcIhZWCh7+
IlcY8in0gI+1Kft3Tv0th0ThcUJNL2rtYgwv2A0FcpY0xmFFm/cETdotTZX+t7kf
OgHCfenQJQ/sMyd199uMQREDgV9JU620tsSBY8W1S/Mlt2BvlqWHTC/nl/vDE002
AWMlsGm1Eggl8SkKqdLg0fYRsNG/twDW2KEVGgNilc8jCvU2hZpa/FaNhiEB5dz1
kjNxygszLoJoxRJ9GXS55xuFWrLIAQLyahpK0ixrw2ryimgzEk+X5GVccwi3X17Z
fREob5Q8uXfYYStG3g7qL82tMviYHYu0S6qiHOWr68pFRJKrhwku8RmT7SQQx2PJ
MbCdH4EJ64GSGalRY4Sc/eQflCuqsXvVmpMMiY5E7bRq1PRgwL3wx4zBfzvRM68K
KGYzDx4qjnrxFo0iGX0q2Lt8PtwzJJ7nZwW9e6/unDtVs3U5Ms4PUX/KPHOTJrMr
B2otKQkzRV50KkcMr6ijUif+FLP9IIpv/LXD0SEhS07iz2HFwzdSaJNiQyKSPuLw
cjNokBLRjJTrIgsZ6jXFhYt/PDamWm2qGbuPp1LhXS8SCdM6oV5XuRHxGdRDT+o6
KH3bSWWhiLtXjuRyKc27h5Mc4lCQ9XydKuttq91ut8YcU5eBXyWhClUzJCQ9Dpiy
gnQmhQSY6EkNOPDx1AxfovH68JyCOxfk4fx3ExPCCJNFB0PCoJ/6OsAtXddbObah
rGSU3XC6rqdTwhqeImJVukFd4fwPLNzukQzwRNfvDtPNZA5QshpDc0Hynn/6aGm/
GC4AeLwTIaNgV3aBhsS224P3WLz+6WJDGde83nibfjVPUVMnjk2jatHqcJTvVWWv
AqGe0KJnju6tjGCewkOrHdbNMy2Nzq9gSVibLNAxHIbf1o75AWVJT6ud+lDZdlTF
0o8GC5K1WabAqjnKICPXJEmHWpViPai9cshpRbhugKw45y6QJQtJYCQkmGLt/DdW
7KmIQmTnCzSkvvpEsdyw1TlJ40DqmhlYfR/XlH71s0avBIDlafZqUMEUeNAdTX4W
KHnxE/dBvNV3ghElgaRO/XF5cn6J9DYLjCEtlR3xvqEHMQw9LG8ZD6dsa/T7coBg
h1BoZT8auiRi4E2OMrYjUNBBL+3+mFiPSyQd5g3XgdxIA77WmWClKgAEMHhgpXKD
T0M9pCqvMJCIVXqpHPr6BHmpB5n8aurp08vFCZrfcFJUeerNM9E1hpWKmWfCYlA1
l0LLsx37HJc0XrqXwTLp+Yh7fjzruXqiX563qX6bLsivxMBNqh1n/TGTguF+a/2j
uCRWApkAvXmSWE7yBmXcQ7nHne2FS1JyHbGHmrlIoooE1VMC6qDqFbb0zb3hJl2c
CndhK1wWAv/JxHQM9UGXC7//YkXF5ZW9PiSQpaAl9+K0lGfDdiPqZprDJqUgk7rx
9xlisc3H4crWR5iTktrcVv/Sj2A++V1iIjullddQkxHHJO2YlShmid2pULl1jIq1
CYc7lklcEDeMG139AoBOCag688pDZQobkTuJTogH0Xfs+189Dm5ci2+ckGi0ZaFb
G26RuJJyJHG8l8GSzaznKpysBMZV6LVUS/vGqFE4sW+YTu869R5cNgzV96h+ut5l
Mf1WEaFbenNIkONJTVSPBIacv8RHAbnxCuBe9UPEpEY+qdnkBEm3ak4suuZ6XJSK
odd1HiVMbSUDHrxVl01/YPNs7fkp7ljOlHqytYmy+fcxRuHZeZKtqotqsglVK8kq
zvIEKFPqu9J4Oc8vx4RJ1aGfrzqYOroQXKcwpaD+HBu1ecXBZPN8hvqZMLWZodz7
PjaNps3cfPbWRoPDFA5voDnUTt4Cy8lCNjPNx23HxCHJszTKjgqICioC1ZIXsZq9
yUENWIhwYix83xzqVBTdEmtzFOeYThHL71aQdRv5XSX683+loW7Cqt534yZXE5eY
mp6qL3iVqQIn5Di1vWqyHUpUVrcaEKTsyAO6/Rdh5KNPrej258oO9YmsF5bI4Lh+
nFo/epLtEzf4GEs+QRww9sbj9StOB+b1TdxGDvdDrochA7ntVGRCta6awUBjevwB
vCt3/K7+LE5Xmn9bZSEh/hsYNygXXuREXzSFNoK/ULFcwAgwalU4iD4yH5NMzae4
DLZWVq5lmpWDWm/i+G+lOSiDt5pZ2b64qSiD6gQEBAFt6SZ+UhL6oQEKUo7uDhrX
DoqSLVT4KWmMw9RlojY6Jpt1xg2oW7ho6T/nu/1Ypt0Bb2JxnD/RM2Gw+wRBghb/
plSjxOTItZS45ZQZKmB77OYVadhyeFUpEfgpKl9opB2iOeDHa3jUrPFrx2wLlLlb
NwCJv8vDzYvA5o2s3esEh2OWfO0SMKiWcUYzgQsTyvpMluXn+5Hn5mJaxxkSBoF8
DtLedsVrBLnYKaN6SgzLWC4QdHT7UibZStq3noexP4kK4baAjk90lk8tYlC1OSvX
5do1lR0iyuTs7RLu596qztJ0x44pQo9ljq9hdQwa+ZELAAvz9/2J7KQaChT5Ssic
Zj0QPZdpQdq3HITXMj3ZkKRDZdTqAQ70ZOYaIrgj2g4w0Gkq5MMDUTIEaOOAvRlW
Oki8Taiuruq5Xlni0l79VU3qwEjF7nHCzOv7n61OQ+afuyrPXZ47nuDp2t27mB8R
Y+pB1639tE8L31FEfnXswqjeVGwQkFzUepDngBeWSAWwVyfzABd+RDvjvU+Bnbmx
S6LgY9f4balsy6cAo33RqcZuXp6082W14znxm/4wQ/1v2gsLn+qJeBl9c0gTdyEY
8oPkzWZFDUya/SE078+0PK7gdHzO7UTVpUkyN2dkB79be2ptX2MZkzCUOBES8WzV
0bn528Wf7DTfs9i0t98OT1sH05nJtON4n7Q/xr5XYV7DR4yr29WUUCtclrqInr1K
yCnv+03cKHChLwGJg8X5pEwKQUqjinR1opN4aQ7FyTIe78LFNC377Sv1Dc3IYsZO
SH1rnfq9N79pt/9ELEED+SC+pRCeTuwb360flu24sngKr+Om6RehwzUtjmAMBFhj
af6b5axgaYaduIqD5hj5ZIvm2EHqU8xbwatK4MXWTnzt4UjcVXSXG8cDV3sVCnQ7
wLMHnPcz4l+VBvX4FRHAAnZxnSzoPDBfKWXxh8fm+/UoXey92jR+mOOQY3cMGbDy
Xe/KGPSCRUn8npkzVRBsp6xN8iiIep0sdtK4P86FbZykN/eN0arqS9VFn5nPMy2e
tbkO/OvTUhGn1nbJfc4yX4ZIb5dHtxWHroYeehU5vAXDivsPfJoBDm13ObNGNqbw
6JleL2jY+wOqft8UuAkeA1JWCFYC+INLf1HCDtA7qyDgML3CnV0QyCQTqlxbJ31T
mA0Wa1bP9mZRr/L1dQ3dB2meWTJRdt5ehnrn3CsLk3KoHujDEC1xZ4I5C95dYGVO
LylCa08F6sG5uinPVm4hXjjETa/KunadX30VdVZ0VH12FAbI4NXXY7h0Tc9KldJc
VzI9NjdwytTC9gMpBoV4X7Sm7VEmX4ZyBCw78oGjhREQjQtOQeXq5JzYiYg6V7kM
fEscLe7MoJBizeziZe9lCOqfvt8og66l6LFSuZRL5wefgJ90lhVlk+D7yd/t98Ct
T+gnwM1r08gEV3xOjuVkO86o21UnKhUslZ3nJye9iXAWGqh448L6PaEJAzTu+G5i
HfBAEo+xEWJECqa4P8nFMEq6zzZqyeSJXOF/PaMqe+ff6fzDlXH74ZpMVbONvAos
WDnwlpzI5bM845MLy0TA2xBfgRNwRt+olxRjhnrSBsg8u0xwUAPPTk+s32rZoW6y
Hsc6SAXNbLsSsCvWPOzOSbymSkZLBl32L5dvZKTDKbmWv6UmMVMpqDzbRg4WM+ft
PnHmUmb6PRc+Qb0IubtCPtdHhCJeTF41QvsFUvwMIxYuQbVgAk859PjkBU7leuZR
FKks+Upk0moNBbEyxd4OODdsTdjMSHtwBwi6HTll+LwaUJLMxwuSnUbbWtfXjJJg
luyBUHg8MNdU4cM7DKoMa7gfMERxN/96ey62/ecVr2sjz3wjBbSm+Uc6Z2++to4R
uhD/HAbvilW2lqPbwDIf5YG5uEal6RKDcTx0EQEWfEU0jBNi/7SNUiMdm0zgSKjj
+Hpfaa65tYGoLZoTTz11hGfOPsM2aCY1w15xO6MJh9Ux0DRbF5fgT/AH72zxDpf4
T8tKuedut08VfkgB4sDYXILsn9JtJ1hUFc6HsPOJg6mW+mdO4K25etzHpc93j9Nh
ZYknpGVsEeueM0KVctK+ZpvPz7r7GHtYLjbjCO3iJ28Rri8qCLXqGqMlQsyQbZZo
EwXY9aF6JiqHBoAK5p+hptWHoUhl/TI3fsYLTKo7ZoTvmCv6ae1zEY3l8nZz09ND
Kz4jVmyFoJXGJRLuigYPck5Jwk8ek7feIxc4qK9RLUDST+63E1LvVzLzwx80Z3QY
pAw9qPISTCx0mTWzkBS4NfpIH8S44Fh20l7i7nE2CtB23kBBe37BYJD85HcL2Aq4
NsPpJ6PNB/50HEzTjOZPJfb3/IURdPUQQ2s5gSH2An7yccB9ALCs4C9apa7lfKnV
0gkGpDOMgIcLP2KSJYcriEHOl/PG8nXcYiztK47/ovzreyFiXgX5DX4r/JzSKcKg
jb+8F1Izfflh1on5Y9dfnkYC3WjMM5oLiH7cq2DQUg6El4/EYl5mEqo3NHE4kcei
QR1oT7tURBXespf8JYMNX58oyXzpe21UJ3SVFR83+gVl/Kk0WADmh/eLJgZsxy6L
mjI9DFE4Yop6bZ6dkYRfIxYK+qtA9T0QwTz9X2ldqpATb0hwPo+aWAGdb9cfYAdk
toX6JPf1VZqucfZKhVbGr5bXh7sPRXPMiOCRfxKDMxR0r8k/ViTSgFE6btM/N+rw
0UDz1NQDyrjUaXKUNP5kjDy//yy6uEdNzDBb0YKCUXsqKPtPrulCxfi518x50hLK
O82+ekG82QHpMqoGz+yTRNyF/STfV3jJzC8QZqkHPh1lkO8/IpsEjN6tcWg5fN1V
FiwUzY2J/1wg2P0QPrwHQ7qhyF4Yl7IIXATaoJL/XtgDtbQXhpqXR5ZIfWV7U2So
BhsYV0Enf+YsIF+xd2Os0ZaFRCXmSrS6KBq74X+xxWm6oblU3hu37jNjuTGMGcGN
Pl2TTydbMwGq5ou+ZYqHnWHveVXThtICzAGqP+rdUnvaNnf9R/PUy/9IgIys1yLg
JRK+iO8h01k1onkblscuEmRlHudiZ0LujfoFYXXddut1E7gMMT8OJ1JeQcgg57Jp
MUm9VnlR8w6R0SmwvQ0IygJBwpDIxRTGUJHkmSnjaT9pwWcoJHoETTLjKnNKBosW
TnlauT/cFfuu0ePwt3etp51cYr74NnUKwiZy/H1klnw/hkrtrr8+xI5w9YdhvYJ7
unclaH17LFIO+FtNPRqTbuiDiW268Gldk38D34BDqY78jAlI11jZMDxi+TyiSXD+
URX2ItKtQt0Hj65yPbQqwdG7fdWRAQGutIsykgakgnIW657Cbe0lsdA4n3zNNXR6
Ds58kAojHYo/2JwJoP01TBA0qpczacnQCDv+s5ScPLb6ZiSkxjww664R8txhzjaw
UuIGHjpc+vGgYVa+1MteVFx9d5Dc7q3tklHhEouSRIR4KSiBGzfdStFYiPDUDMwo
l5rgPZCeNIVW6zt7Ph4anE5uc09t6X/Ej2KaDEHtRvGIsBvJ3mFFx0EC9d5maUuE
S4eOmlPy9RGg1E3MB4aAMOEgsdnBMtc7Axb6C3i0H22jJGM5POfdyxYCSg5dfvRv
SnuUQGydxqw1mw07uEOQjDhbc+qi5J/3cN77EEGsA+rhiE24Idu8JGktgZ5ppeYH
zwYyO+s3kOSjjf7ePePvRSNpJ0Zc8nH9f0x9iRlwFL3dRAzZ89dh51vyZi/0l8lk
5mIUWdQ4weXzU8oRtTC/TjnNc5PMxliDa4aSuSS1WSzyvKqCqJA8onbn1/INtxNM
GcDRfzM/S7+TlgcIgzBe1HOGJ4/BPqBKqmNRypNbY0Pvx4yGJkI5fv3Y3BWzo86F
CHdF+L2lbcx40SKKs5DcUerMCZRJmkuYICv+6aApBGSaftoBKCJ7yx/e/cuqNYl3
f3Toy0f77+MA5vJrPP1j+RZwGiBMKxcJE4f/IkvrZpdJTM8bJumP8rYdj8jpXGoO
S+w3f0P+M4ELBN57e5tBUawyzsD7DcJ8z89BZ63BKbYilhz7qcugDdCJxq6QxRFV
AFrfJYlsnmmTFSGDgNMsJ+MzkSFJw5y8if+zbKjgcm+697dn1uhO+5/Rfcn009Iz
DMcOOBwB0c60Oh2Sj2d6YZSNOg3r0o69heczcuZl2ews7EPwJmN+jbEtogfeHpKs
8UxcHQRA5XHPVxBUuMDW0z0MIO8oIK1QzPOfLJRHPY5BMrncPZEb5fo/My/DP4bj
ZD8bhZDDu7nJIMR/3wyZn7W8LMQNdqAtK0416aRkC3S7cyzwHKp7bKMqewHPOcxb
7wQOx7tMd9ONaBBhHkXRo6anbqxNA+RdAjz3651wEAkj4qgNUdqYyGPSYxEFn2jQ
lF4Z+zLqOMS3FmPEc95GUFT0pIW16JCNMtpWwMsx6xmpxxnU0uik00iTHEJ3lMRI
1MwBdt+tPwBeeB8d2FOPDR2dlP7oMhn/76ykFA76GNGBOJqM7WnrkFT8TKjvEXuZ
KjbdFyIcZ6XBguXfQBrsmGRSXViZWur/17wrvamICKNcfxm2DWjdGtYzuvlNrhT/
rveA6zQd2SuwTpmJnYvLhFghEtqyoOrInQjYDbphC1T7MuuIKQTlcwnHd9Mqevd+
WDt+sAbRfGHmGicvg2j/6vi6ZecV92whEcuF0PSjjSDw0ZMiwtNMb0cMlZvOBi3m
g5QXm+j6NJc5hfEX0dViUwKgAWE4g1lUrlEUYoKaIvyehjprxch23+lWHa67IuMj
rr73XS4eeukFo8/1IXJARaCfs0nEI78zpPRyqeThWBb0OXo/ZRnewWVsiP+Hi3rM
ikbA9U9ECmulh64SSrBquxU4nAs6ZXxxFlql2cYVGxlZp1PmRUSG8bfCu0aBJYxh
iuaSdqjuj1E+FTbru3iyni87o+ZvWqfjr2erntbPxYMlMl0TFPmT3lpfl+pa9pm9
pHpaan2jBu2UL4e2EVFvz1KGm9uxliFxvCmFa5F7DiwaGUpS3M7XDV8+oHSqjSGT
Jo1raIF8Bv1ND6+XHu2OAYOznOsVkC8KpnL+b0xNwml4C9PbtzZyWOkdptohovGi
RcuSj+e+TD8Rgsuv8d77LU+QLvDJL5lHRANr+950wXL4hdfMAEFU1agQxU5Y1zBm
LgtLuQfbYRoQ9Fh8eXEsgX8CHntPqUMKH2MFiBR+kH+wB8CCYdHd6/gVb86QhIwv
BV1HG94WRrpNZBGozOzoX0ijeqGmSgf7EglD/4clkt3DOlohVmTgCz5e39vEm7cF
X5oiHZLC0LFXvfaaQ9rcLjAWjM6Vw1+3SzrWQKug3Xr1vMnp0/tpZItavAQ9fofx
+UY3G0AGEb9JGobBRaQz1gbiL7MsD04xsjNi1/b4vbJA9/rUKo1cHuP6hIwDG8Co
Ujy+Kkl0UO1cs9IP3CQvTbHgn1DWdRoVadBDcJJ/zxSAvgL/Ax/6Y0LfRqzY1EWx
+DkIo01w9J6KuogM6Yv00vod8b5rijMDQMT/NAiX7W+lqAyFPWBTLrRp4mgXUMNi
AyAVXbFSy4VkbcDG73VcNPR9nJOz2zkd2uWuwoFtImAri7GCH8N6YpqPV/mGVOwn
XvlRJJHDYYsXPCiBU2TMJ9Stxwgp+Tn3aU+Cdd6PFiHgPVPwyP0i9ZE+Mt/UgroD
yhzr9uruuIHlgnUv/ETnDMtc6K2NCHgxKaiqu2VDujMyC9qJQhFyap8fumH4CA+t
J19bAoJYqEuinwE5AjhGXp9wxqI4SQqPN0i4fh73XIX+zJ/eDzfxZzfYhsaXmiFp
745Nk1u0mOc7evSpq4C8dt5ZEAXV4Tece9+RDBuB3TKpL9pQanUPKVoOQf1x/tzA
uU+x3kdBil6COwhmhCIWo9J7Yfan+41FDFGOLBelvZvFVuMLxGISPBj9IrpNLwjq
VWLhGYPCD7mfBTy/YE5QdPKSRYkCcyT7Svf44e9rAdKRKA9iHbDryixZdayToLQK
vmACl2CUhneSvIFfvenjMbHO6DlxubL1ACB9zTuveN7sg5IUApltmBsMHoptNAdO
QsOpEsPJmjJvO/8tCMnywXnn9qkRZ809z/U24lHGsPGYo/Nu0fEOIUje+UAaHfxO
mQ+S7LN59DibAJFhPW3KIP9zHMvgsH1OeE+9SWoggfp8PnFYhEq5CbdhStHNacj/
CazerfKOQFfn/385XWpjFbtkZw0Bf2f6BbH03u9JLnrWC8z7gYRcomUyRWYrlk0X
SuyfWxnanSAyZizPFyzqGuhtqh6bQ7PHx6kYgHmkKicHqdxmPJDqAsaizRQS/CMQ
heZz37UJvw06r9FZY+bSB8KHYnHedQmuuoFBlpLIF1nM6/8LSd4kXnF2n0Ek9Zlr
CcnGkyGYmd+0hvsj6oYAzeBx0blHAy9LHIAHYu27qx9L98SUnnLeLz8zIf/2hF14
8f7Wz3cvTBuw4FqnRykr0Y+BttmXgdEORHT06GLQEuoQrImvc2la1NwXFduxp8jg
TBMbLwVczK4wry1MFK5PvhTXYbAcgc5qMFPbs3ql94fEGXjjwjqLe7XLMQIOEnoD
ExCzlZrESBXDfA2k4pf8+jrfFpwi3GGQ/LkJ+l9G8uHTJeSQKkvX++p7lKUYlwwX
XETG1L/XMnXPKHgCi0k4c63YjQhQeM35YdfEffT1PHkxmeE/NQPjsMgDm74IS7zC
NwFecrBkYS4/as+mjt44JYkpitUjziv4UIRZr/BVaT5EQRinISr1nZkhnWWH2Ocm
L0oRd3z4ShzomJl4aa3z9r58Wk3LcJyAdBZA8PvQB81IQw5nGe9jrQKbfEIAcPr2
HjRjMT8201yL8Di/CEj6HqGdDCOzwQwmz8wHsxt+x6IMmD3xqa6uaaO0G2NVkjIc
UoRLoSk87rfpdWvzBLhBe3T4v+byIYmA7ZscVxa8/QJPhA72ECbI829fzJz2JWMt
/L9d8BRt3KjErfnKRXOJ+3XbfN9fCw6QC6BxISNyuXyE6/EUQCs8WMQCaZWWqwbV
/30LmSzac5uP8T/U3Pw0ummJM0NS7XH/JHCRLV+Si7vi7DxUIEzV4rUjZSoXA6ab
sJeirq8VWBgA7qADL/ByGMlwYhFblnBhBrRdVIPlO/VU8HcePNPYiPfaZf8Ef/vY
vHvMoOibP/9uRMAs8gH1wPn0nej7tevhC02aiZKFdL5NkdZntw2eUD+c4qKewLb7
4gkAq3KIpJ+tk7QA5kqf2kmQvxfIWa0XdWmAelBzxbIL9dKrsJ3YtRtu1BG7YdUc
X2LWKEdlfbHE8VZcimsTGrmh9zd0+I8yBrGnfT2CNUkRcv5t1Phi6DoRd8I/Vne/
ME39vaSq15QPm1TjC7EjiDvF//t0jB6dAhuYVmYajuyBcFHor9Ezhjk7AL8lZNl+
bjxho3kLTiqGuhSTr2g9fLrBOB2JkXkpJTLUb8RV2BIjYCXO2/N76sOVn22ckakm
EZ91tliSycKtDc7AdftBmn5OxBdCE+k+G1YgSCulcBEU52OPkVG0aveyaL6ba8Br
dNm0K6ScEmNuSfDmmkNuuTW9rmLb5tlpA3IQi8gQf+mBX21KeLd/JnCUXsjyCFtf
ArCt3ZG1+a8EWJWyndCJbQIIkoQs/X4VH1XGMzOyL+lSRAdXcHtEski5t4pFn4ke
4UzbJnzoKIjct066b/ATmx2fNdv8D36B7/tWu26T6ApBedseo+mba0NhAV6ZmbSP
HohdmkUTfDpNdGN1h4x1p5uVaLk3GGPxPwYYPdhX1xId7MLzDWQPOwDBDPjxgop/
VXo2l7/jrP3nm/i1i6f+ZY6w/eoVXeA2hUmUXVinxqFAlXd/MkxFE/WSSJncxpv7
xEk9X2bp7L2nhJKZlyP9lqoE6tnll6CG4gIlxUMYiv5T9n9xSWcN029FqnHrOfXd
hhVY6a/O3Fh/KmBQ1Kcpe0bkVpJGtQStGyc66akjdT/cqK9nBfd9d3Yp9adIvhBI
KQtOhoEURiktMPp6ljYce/HGF/3pCwaTlxmOq3sm8N9yXff11hLVqyAmqNeSWKYF
UMNT8ab3mQPehMczdu8OsVOwRdAh2sXhck7eXd3UcfDUf0O/7mSub5e5yS9qtf4l
oRRzJKZrREFUg6SApH3DCPTW9OshvGS8mqWf3Qsgr1GpZo5rOg5y3Wmv0BG90fT1
uLDlrYxBCD1KFOQimuot5e7Fwnajs3rR3UdkTAVQdS5DBxpKKyvyyTauEDm25vQt
MGx75HARNdCfUJ2OTCLN3nu8XGxWMp6AZk+fvKoGuaq+CRlPTQHhXkL9cX53Qa+X
Wkt5pSHMyKJzaNeSR3pMnQfWNu1/A5usF/YdeFupVuYm1RpNYi8pI3MJc026hi4+
11BctU9Q+Yn1cMeXWv51Jqg2dVI1sqzE3xxJDl45cb/qOEzXMPGZ+NDGkF+dB+gh
kjTZlDtPaCbJb7uWE1wMeug4b0mYGLdRtUJUjuJsTmnFbSRNhvbD8HvGPYP/h6kX
0d7mfKCuvbkj905IvimS7VHz5/B9ojIv8IaTRl29N6G4tmdLttF1JJ/WE6dWERxd
PX6wTE7e0VuxiLdfGA0maENL9GpVKq19eHGm4Y6bKHyUCZ59QoKNyWNZpXSf3YiG
xOHl5Kj7kikzrWkbL36UJpT7oly/EKEqJLKql6fJWPeHODXnZ7Rk94QS+jJt8Qok
vStzU6ZcZHXUpY0lGCDyi8OJkAhZbm1RXOlAkWPzQYmD+p7Zx6nZ9Epy3ubMRTfR
3kTs62uCWy72OgIgF0EeIzMNcNhfa8EDWopkzfsIBuM5pSzIRAygFwWUHIAqSARw
FYwxA0DQNtR/8gogyA9K5m/sqVdvR1l+/3UpzXt9+JH/btBNfSt7UhxiJLej+xVk
XqSyOBO1StlTYUqXOXLiRkp9kf8i52goxNsor2ZBQNMyBGtDeRP3edQkpFRTpNzM
2YjbI0eZFKrlWT0weHNQsD+dZKD+lXtd+XXxLWRke4vsTjZZ+K2t14Ypj99uQs6w
zzGelzxhe55k4eD/N31Xv3TZUIgdRwadYTI/GiJ6S7eNM/hiUOuxHa3qySdM+NGW
2F5eWl/NBaEAQtp4gAjEayDYUU+XiCF1IZNdCUh5AKYd+tHmtnoU6emYT83VYXl5
oJ0h2TkImxp4IqPhP1GJXUra5NCTuBAiDDCQfp/svBUCMV7wFSizNHKrTHo/xseu
aPae8jejJrKvtx/TAE70axIOS/S5JwNz+qtmf87Y1jKrQ9OVQH1ZP76anrx6iq+Z
w7pQXnqVqg1BNJYbrS88lNPaT7w5CpTLJA9K6KfPitbXKb6j9RynnftcZcY+JLnV
SnDOAD7a7Ll3aN/mpgdclkW/d8BgLfF7/9wQ9KOypkOrnhAybex4VmNhkTJhehRk
IMNw30J1KJNXywmpCpFiAkjQkdYlnFNHa2ualwOmjihZn3KXaP9A5tAx0ehYu+KS
/bawIhZifH/2v+1EnbIbc2hXOrugCPmclQ1ATxxr4z73N7IDFSBN7Gk67qhb630f
7SmUodCEk6EjVqMq1MFIO8A+APhZZGfW8vl+CG4GGO6esl3w6lqeW5Blx0vpOxgH
f994CZlM3SCVvEGSTI73q3FaFWKNdoobvOOoNEYR/Gw2sUK9r2GFIhACCQLGbU3U
E+mqEzwOauiJSODa72aGfImkGUiR9vLu1FW3eUaYdKHqIDn2xZnKsbLXt+PsvL/h
km7ewtRg3FF0UU0ReBigG4p9UaVkDo5eRSL+KilkUbIoratgIZRusxdmSOPp4fIY
2FI2dVPdRFVL/hFbJA9MuOuuMus9eAWdm6GUrr1twWIirt+tZEoNIDScxRWQ9MJi
xqkSN3vNf4795Ji4QgRCJIdKnvaCglGCktJlJIJOpu/6qScrIQIL6rdPzzncbXYj
H55x9vVS2S4unP4l7kQBB/EhrN5M2SdTkETgcojlJEM7tfxZSyCV7VZfeR7GE1Tc
6w0ODeUJk3EBAuoBKH93H2z+P6mRQ3Bk3Yn8YT6NiMqSH8N1vxGpRBwnAuQdPFF4
Z7JF4mGky8ws6+NAiVSMmofW3HK7gMM/ODJ7M21+dZbijOkv1xqSB+6JH6fthmIV
3KVzor4qGezIGD/fDGEt1ovB23kGakEsGpOc7/ZmfigPA+65anWn9lxAvywSPjhg
AaXthdCwvTM14tyohdgGMpDEzBH7qWJ/oOMqJeC5GT/bHVnHn0/w0ABswqO3oTNi
BTEFaWmH8l3yw+EfW1KiLQarcB00kM2G5Pc2mFYeA6f7KHvwv+D4+h8YJj2DJ3YO
njlj0sCJfiaXgYBRZQGXblzXGKAgnGelJPJ47eTXvsWVOTRTnAXQ1NjLIqqFQOi0
p3313edT+MAwJ0zhZefgJ1l9xeh0crpvp3sNvMjDoPP9OusdK0VVmCNl9YsGPr5F
dfCztlixpKulqjoecBMvqGjURXcWfdMwsD9mGJeF94WOnF9uYMakGp1WtUoDhqq+
rlUbwFwwoDUwDu5+MJLGH3xbtCMtvYOlIVN9Qi0Ffuf1ZeoDLjtIHWeJGucIpFsh
DK/7+u4yXmvbGkWZze6kMCkadYuCXXgBjLK9eGc394VRYgmEMkxo1/9dmymGzEmN
I7ft+Kj7OTDAWzhsgQlttweCFmumLQ2VQg6XH8pEWtL+J2wEH9sAKBuQlBd3CdQb
MTR1/rKwwL81dLaXK4Pil8fTAtoaB/ZX1IqiLeB5I95JZ86exMmSvIUzymjN3a9N
GLBiNGyxt2+/32gJm5q4G9F7wHc6Be9+Y+6I6u0F2r5n4VNatyfEeVHmv1rhdu/m
Jqr5LHSWBRmyZQ0cHjSFsquyJO2VBeb079vDl+FshmfEbubrgqhQBSuVCETVIVyz
in8N84BkzqrVqdrA2SVCP97QREuHUcJ9l8VFD7yzZ0+tUpFE3szA4qh/DDT2jA2k
YeMSv0JUA54Q2a5dxI2FG1pcerGQ+NuVUTQsyV0pYhJ6pGPukBTA/+w7ehRjeckO
tMqy1o9LDHQ4fLzUu69KnWH7l/iYgRLuJz+Wi09Da6VJfUUAVPKoxFctT0+S2KvR
6nSbVSn/YMKlBJx2KoNKPiBcaj9MwFW6CEvO+r0VYTr16yfVgFYwXKdyx90MbK5z
eovXSAIdLKMdvcUW2LVMuORelos4LE1Z2uDeF0JjEyd4Hi+3oa4IPY126MARmZb5
OZBhXLIkHGsVq6zY8A1u/P9MxZDU5eUvAxviEbPFCsT989nQn0q1qvQeaMMiRH4c
G0HAmzstisYv0JUlH6dpiTCF/tzSp5ziXlQphoIgXGHhhNkQvKkvnWW6rAZfTBr1
wRQkoSehDLtJ28oNzWsAHuu4qbokn2OvyMkHAxQQSoXQnyisqvJcy7k1cVY9AGjZ
B6E/yhykSMmAFFnQOF0F0oMt+DWgij+S7EoKXIWmRw9xoOO4gM8+WLuKlloQyuCk
qXn16pZ660RbHpOUm1sYRGMpW5OYnaPRVbzMZ41wHJ8uvEnjzp4gNMZlD++0o6TY
clnN+2dDzNxZ2Yji+jC2QHPnaV6CW881by6kGrCNYGPDbH8EpvFt8i/lbIwJXmvB
untE9Ug/24BbLx10iT6YL+eYCotbhOKKssfbSVkqfFG/AvOZH2AmyI2rXmM4x+b9
OG+2BE7OqM4XyBezZtiUigY0eUe5u4uNudfKPZGNavSQWE45bIaCA30IBZThGiC9
wgALx5H8jIIFdV+KQA9NyrXTnaU0un0o44FpvY3q2hmZGM+b+r9e4o66+CRHwSnq
xhhIWA1nQ8bqry+FOc8NM4v+TpS8Skqfm1bBllL2F7KEQ7Sf1QpXPRFDQh6FZnUH
2xuam7XMGudV2CJAmQB+PsH/S3X35vkjH1wYdqy6FCjVBF1UNRqGTh//IriPd3vX
QEWBo3nWjQMMdpI9eSBBXTCr7dWtevcgtQjxItWfnOxDyYJjAGExOJmvKYbsRJ7T
vku/ph8xDrVCkmSYWKaYuNPQD4B2JdIedxaN9o6oICNFt4qduEi24HFUbbCLwLsw
pFgw1Hxuym647dGks8nhCJVGuFj4mcMekPRwFHgVWzzl7vrLLqZHTG3n+Ukz2LGO
LjKakDI6s1Ge36xZWlSD+XAsqtWgvcfs2zGJK3NkEcNc2Zmr6X9L3xuLYa6nF4VU
TQFbLV69jRdw3jDNTB//684RvuZcGK9t7tbPxJxcLFc+hd2XQ6WKLoDooSRNKsO1
yFAsk1gEElj3fITK91H3btu4qiIgp7ZkuyTVYfbW7eQDyFdYw1/WRL2XAWrdQjHg
oN/FX/36kR5FC7uP/VbL3VzKuJgG6/qRtvQ52Uv2Cr8OIEh7Ue5O9M9/zxBFHCC8
4kOPFvIFXItG/YyXUmYHoCwYUwIWcXpFM5MfdXcSDKaxzHrwBqF/UeViZGtK/xbS
/fE5D+0nSpG07SsiweRp+rE4l00cg7mzXTXIZv9ANsqOHZiPLxem+Ks6wsOznQbq
5naXJ+mOAxJGRIyt0SHyQnSBKQmVd1tIpAhfXAjIlVCVE8ccQOasecoYMFuz4epl
OyCvKYXn4kOcbQe1KV6icmJllcjLj6fM9IzeRy33FJkQiOqT9zaUgM9P1MKvjnq8
gh2GndZgzgPy707W97PRzSwyv+f3skUtbolPlqnjzPkr1JylOyJA5kJiHbtWPKhJ
t/TCd/dqeic3z5qbZq6pHahHUIcpONTyeOHFrPO0KH/vbONl8IcahaKaSy2qpTpK
PLWHgrvAmAJE8LJLDoZXYHnbayjM9tAW9MvlyRw18poDOC9OFPDud0LjNpX/2aV+
MiZLoHiQXxpKsr777VoQdhmRfJhwnL9eyQxVXjsbMLK+wqg1IlaAEI2DJBDF+46w
62NrudL97JP66s4YRSCksp/OZLFFtkjpBtztN3IAludGXTCpo8p60fpCIX9SZurU
q//xPKiBeTE5m7dWu5uiCbeqBr8LSepnQrliJqoSBt2dJ6KH1JLsIiTFCqFpLaNK
+4+TFw1ahy8VfZAc7dLZVOzQE/1fnyuTTSQvuuACu2z5TQum0RVxH4BEha9vi50M
+lEBcvDLdlJQIp2LRhOEHAxVU50ZbjybCxyrBJ0qX+DazMj32XlPWRoJyyEiCaaa
wO4Xgrka327AWkvF0Yf27lKu3kOlh6OKxvStfGdzHqyutPdrbAzyombh4QwwwYoE
4JPnCAIuvSoju6RXVaUaGOaxFy8ppMQS0cwMZ+HmnpY5m/xFxH05nUFZvBH5L33R
nSBZum93AUyHJ5qYealJF0B+WC6V+G2ybUCLLN6LkvRcNMZVkM5W6RHDHJGVBUUY
e/9HUsvOvSBC83q9ozrrLdLLjkG3KS4oAimyJ3Vwej0k3mc2PMh9kQtnMq66agT6
9byK41UF+9YhTwMPTA0l3luQFdu0B/NyIp87uAp8xOExgGi8YBktJvmGxM+KbggY
EnRadH2lU34R/sKinT0naW6V7aIn+wePevff9PWjvxtYi3cgbl5Zy12spZ1QtcH/
VhnjuCCXOE/LQ0/1M25lPL/WhlHN6Xes5FIqbmf+snqInp2uykgECekIgpA1sfhT
j/VTJ3o7fVV7KVwu+O2xDENHInZHOrjrmd9eKM1rEXjYmZGMHrnanXAXNQJer9IC
/xLsMy26r6CfI5Amjuqxx2NkiWx2AHB9D7Zq4Numy+uDzxn/f+mPu0GjuLtxg9Os
uW6NZ6K+dFBw5GuqqKy1r74QWfJYyas17XfS/iSVWj3RLFdS5Pz0ZYZqD6MV2GXw
IdIMMOgZR+sI7RwxIP7k55mU+Bmsk81TWllB4XdaNZBx/usFQlnGpDue2POXt4IA
6X5stJk3mQg9UJMZSe3v2/AkKRd8Jv5jXnfTpeMBv/UsbaSHRjXSstcgcVD8xjjW
VzdSSU+kACJmovckIlxeq5ZP4XGkRFA2zXJHhB7NIR8r+AFfZWXEOFMIEL4XbAjS
R+V2TfZ0ZJW5tRqh5/WrLwI1ePTadfH8OO2pCy9nWTgFu4804tGW+SqMdw7SZVdF
8LAU2VXN3LoXlboGwwCymFDJrhZ1jU10J2dc2gT+/MYSRRVI+xT5H8CVrHv/jXAg
hfsTKrUGAv4OnCkB5L7z9FcC5nUY4lbSNtbpUWrsGCel1qi76WDMAdq1YwgOZMhZ
HNIWbk96gX8Xg8r0nGE4/rh3WZJdeowaMVSPT+UqihUhcpGRI1+9OuZy24VHbuFT
Xk4z5xZ80xxIYtht1pKMaNHM3mAs88jPNyH6tKAqSSmjDoFDvoiWF5XgAkvCZIy0
/j5x3TkIRHCyIn9bQggVG/iWAp31H3RFa/BdmxppyNP/ORtGq/lWUiRwcVd5CUP+
S9DXY06PF/0V/WH5jPBK+0envslZZbqQwVRYO3ps6uF7ebZDYLIGbc4/R2obry+X
s0TJWej3WR29xx0ClWs2R0+a20wwmM078ruyS2yG/kQymx5iNoHNzNQbNOMz2EHO
W7QF1URmN0tb4e5N32oMGOkdR/gdqzEnuivU4J1cbNy5qA9Xcu1xCzgJGQONbUzN
V0TaM/g5vZZFNXPBRykyHBwSQ+7fj6VdiT9n8fNe0Oh+gHSJ9zYTL0HM/FIEmZdH
FgJGgV1n11544xrJrp/RxAI7RgqfpstgHG8ld5QGSkMHFX6YreJCGCpbOU2/Gxui
zsegcckJgKpULMnuFJvV4js0mtSzAgdK8OmWdRueZY7i4mUTlQsge0n9Y8zGIhOi
XoJUrKl8RszHt6417e5ZUSTET7L6beVeBR/+6WWHvYspdez/iIcQ19XscKxxPCru
O6qFbw4t1KimIIQjJaUmQ0VijD2VSWKqf6RnqZInR7PaHHSgQ+aWMwrQCOWDpxHb
3T4smc/IDfyGQx7GLFVX1hurEUCBJJUXZP2D29kvr32ceQmY1ZXMKR9c/46Uls39
HNqEVKavUxtRA2JTwrkpI64rBXVydY2DK6EqA5BKXOpxRcfun1fsK8IFqsbaZpzQ
YGBobi7vpZCPaOrE6smBSK/85GzScScdFdxA+SzmY5fbKYOIb3vopkVEwyfl+GbA
kdx/FNpCyp+JaGJjGbqXEMW7odpMu3fAtF2hmwRLIpOcXQQgTV+o/qPgRf9BijjZ
MxaKfxzbcF2i6MTcYFI6VM2kO0/vCglB5Ni3oHHxVc92SSZ8z10J5gKcKnQoHqU7
GGj2cBwHrfO/EopbcY9MYbfDXZiVoKHNXjavpcFlGWY+rvs7VV8U3mn+Gxn+/bSj
rvS/Vk8X2nAPxaRfRBuzEFn12FRbciXOSOtilCMOAaRRTCERhwg1qn74AFsWoHOz
LxMRGaqsGT0tGe5P7y3FSET8Mzv3op5yIb8eUjiV+SYp285Q8Jf8BeWbAZrWrGag
3CyQREoUDq4DWdWJ8BDby+fML02VO1wbScFkEqb4etYs3Pl2Z/6+v2yds9+1k8DA
1+1EV2fPF2VJs2RHqEs3CFAUezCckt27PBzYqXw8PpbBcjaRQpknpkYJipQTmh+a
lZXE+PHhygJTs7zlqlG/sWuSkUtm94Ar3h7Ieo+Fo7mmdSQRoKodzi8p7ZSf64zg
LdB2SS0Fcglf5UJPJgoU9ZlXJ2IhiSlzdjtdlefd9cLFjryB4KuMwE20IutwEzAi
LlJpHs7QWe5akrlsJeMoW8scV/tOszJ/3Xgy/RpshWLQnl94cB5VAEVcRIaQvaT9
tnAY6kG9xObKR427r9Yw9aL9arg4A+1a+crgaHCCwHhudp0SFBQlG7FfMYn1NalH
MoyGwGKj3jH0OuxnRCNaftTrswUoMJIVf6bw03x2m6Sg63V/s0PfayjN7MRdTDQ6
R396B4z9Iwbv0qfzVR487kTIdczyrFjUr1uBaVjT8DHpNafVMgHDIxIJ0oUG/69V
hjSLd9FMZpokzYm8IofRwWJVVqGGJTzD+CoY1rvIgq2wucXCXLa2tpW2UEHjPd1V
+XqxHJJkUJLqGvkPN1ktl1AHYAxH/qoDIWlzrcYSgljASdNJWmO0ybXs9w/+eC5o
k8VISvrCLfaK9OlBpPvFDPIhzcgu9RSWHw3bcB0PSuBLkKuyNQwKVdF9A+NG/aJz
XCkE0XLINQJ0d0867ty2v1wAdITZK+qHZiDucRc28Yz+z8q8eW6Ao2mlM7qjHmKf
JU8Y4afbkM5Vnfp7j4q8AJoIGwOaiSkn598KbyUpN3ypxP/CvgS1bP3oX4hN34H4
tIN5cPaQGZiQrKCafY6KTQhhSbrzYdTLLXU3Bn50y+jvDky1rF6gyflYWwUnIxGt
etWJ9Ln+swPZeUO5XDb1aI/OmOTvwhdPBSkEVlCaZEIylktOaXC/yq9dYigXADBF
hkImqpcTxKNTQJSS1r3eIpYDuk1nY+fYtW2jx2DAdidp1+4ThawFEEdbwUXkv0ZE
AUuiHvUZaBC7dUwpxA1UaHwJPR2bDZuX99gbSVN/Vrvn/yHUjn43fZKh8LHxZEhA
X1F/4koPZQsHB+fqtc0/FyIvOR8rrHqzqQwSflvFjkYcvCCehYPvBYD3XQBeybWS
AkffIjN2XDk2QX4V3/naHaX8afEw0c18E7NsHMBBFbTrNZyKfh20WhD5Q7+k2Ral
6SYc89UgR1YcL4crL7AAbAGRjo29zrqq80dqdhzihCmOKpAEf8649RDIMZWVOFcS
xwqUYFsjaZG2WE3qwhlMG0/beSJu73shpjlU2gv69pzfXdEE7uTf8Taf2o3NAj/c
TMKRNuWVja1PQ0w44Tj6+koO0QPqrdj9p9N2dG9liaIXY+PHQ95VDBc2AxIVjLjq
zdVrEvVufQCqYJhEuNAjz3LROeCVJBeUPQ+ZpD1hX1bbLdmEvjPZwqG7uR6YU0NF
3qHcdkEw2d85gUmSFaUYXuU7BpTiNX0X4H30hrNArMdERtWqYr3AWE+hfzXtpCJg
p3md/1uqCfX2YlF2JCiMsoW2FjX/02vFOxmSa6kx/U0CRuMYZK4wLiFqsf8Dhgt6
j4EEQWvkib1kYKpgbERcjtHo1QcETXria5KDKstBeOhGUnzBbWoBKloIHngrFVku
o2bQvSCWxzaCvmJ3ROoTpnelRcsyevwlE/DbQ+JiS4YycAOwwkzvOaV4WklGT8om
m8eCPUssDYz+7RPdTV6TjBUV5XDV2quYPeh6U4w+jmz6EIHYqp9BuwR1rA/dqUUb
ZM0dTz3NoJef6mSVPN5ENjSKKhKSu2jCcYk0mwvj9V3oAIl22UM6VAj8b8vpjMsQ
zNfF0J02jitfa3q/7vkc8DLwZu0Ww57J6dbW4MRldU8MyDQH/BEoe5scWKlwRgXR
LFnffR1xI+904RKCeESMIdJu/FRqSOWn0kM82j8Fjd9PuGQDH//lKUca2JB+B63q
9WdXgLpOZxAYbzKki6xlOLtqmUtuWKaZQhgWj8rDi6iYTqV+KW3yt1npcE9dI1Lu
471rGx233NP1KScI1LwbDwMv91T+dX3ZFXF+EvF3Akxj0EVqeEVJyNDLwXbsLLQ+
+MVvX1Cd/y0LGVxBk6uLKyBiKdh+TznVAa5AKKiaOfL/z2xjph9fPJmtwBvV90N3
hry0DEFkY1lSVRMsHUeCpBZ5yzoHHKr9dEGseKhUDyu+tB6hp5UiYsdYihP9jXBj
7ei3kzOCixI62qbq2712GbNO0wF02KdBzNMAYqE2qVEuwIiKle/Vfhc9irjltlDN
jktsRHjBQotpAS+6Gj7DScMUm0GMfcUs5ghrQY4lqr7kkCmBXgtp4ESxDEVaccrv
OBOH/EOOnsRw9QkTVi0JposJExzHkd8+7qhkYFNl1tYigPQ8OtPeW10H8jELnazm
kh91CpmMsjQYINlkLRhrifLpwBGA64wVXIcNGZ4BEbU+TEa2wDe0R0tQDZ37qnFj
zHYMLGwznsy8dzarp3/smcmd0iNi3/KqJ+aGSkYt7NiRDkG+Xbkd9buTYTmkfUuy
+OgLeJOTiURlmFJN66gr8eotMW8hUBnUC4uN0BFraTwS+hCJ2xGmjGlorRNknSx5
UI7OgOC5pGA4PPD73IjwmH9a6I3A4G941TW+797Y3gjH5lBj9AA673QCndSZ6NR+
vG6ug3OxLSdGUWnclmH6G8NJexCt3b5j9EoOzb4o6/BufB6/EwElMAnui2KvO0zp
jGprOUN6h7A0Xbk6ojaiSDYYSgHQ+n64ykPNPuHPA9p2k+MsYWMbxm1SBHwgBjku
S4OTqA5uMy9luRD9fUmI2Rk3XI9CbxirJ5a0Oma8mXRGpylIMmUCWuCvsANow/ih
SCNP3s+mfe0lN60CCHsOPpNMNxzB9L5bS5lAqcizbYhaG9y85w04azyNq8dcWvgY
XDe/R8aKg3/JBlYjZIx5SDOijyfas1ONG+FIzSVFAxg+bnNIPVxpYjqyYXCyyG4i
9gPuMyoayY0xoHtlDN7mjfAtVJgdrSnlN7Re4YtHWduVSWPzCKgVaLHzhUjprPCs
DKtRVJ37QltSBK1vnTRVDkZsIo2aQh4yxoCh4uRyt50Vacxcq2ZC5/oyFFHK2AiD
aK1YxdGUdzLvwMB1SuPcSc8ewe9c/clUNdS+WR+6kl+n8yXn+ci6ZSXk+PAq4jLY
+PQdhFm2M8EXzEV5i2/JnkvVJaLhb08p8CabYTyUhDgWW8/BWdiTn8rknwKIXNwW
MJ2doEVxaE3rwBDCHqXtLl8/FbqAYgnDSJKCrKpb/Fk3cG/meqWA2B0S4CDFLqig
KS7BTauBuABIoFkMaZxyGSkJAnKb9vKrSb2Yp5JiTQ3IRUNetd1JJIY/ZuJh3HWo
u+sTY5uMvQ1qVW9fNlJPU2c2j8FWpUs4dhZPCCktm/UIK0jgH3zPjYJYShOOXNP1
FGIArmZ9UGrs1esXQeEBHA2x7kClEWNw4wqyJFBDY1USnETTM0MlR2MOv18XL7g/
hISFU17B+RrRnxqiOrP+BKSLgNqHqD2CG3vx67x2eh3YvWud0RNNVbIvuU8/l7wY
Cvn682tNqtzThHwd4VTi0G4cFjK43CBhfD7GY53DhDGdECFMNZLiPIVCmCwnbfy4
8eK6WAd4ZI8nVdX3ad8UvlDUASqCMcp8FCAUtqGd+WtzweRCYcuZcCcQqwPCxHzL
NVMeihjWMiYpvSnDwxlWlYQ/rNfjXEOj3j82HNmg9aST2ayhxG6WXgEVkk5JxnOT
Wda4WIuWaqVgGgMD5RhuVlYzK0sxh8+a9LN2hQjJaIQHOrvICuRi173S6BMReWdj
msutb1aeg+KRPXSa/WsjpshRdH3cwHk1fhyVpe2FOj0itftE9slUFk82rGp21ek1
HnFX438qK1qpPwQzdBM45VsuAX/FFlvV77EpEmRouWk=
//pragma protect end_data_block
//pragma protect digest_block
yxlf57t+fffXcIPySbRSebtC7Mg=
//pragma protect end_digest_block
//pragma protect end_protected
