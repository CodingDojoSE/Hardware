// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
L4lqMn2BM3aHZt7VwwGv2GAqd9l3l9ELZ6AeGMCm2HJPyPgfkeGv3RhjehE6hZGGHmnE+DMvtwx0
JSrKzRuXq7WKiPU7Rz1jywkBUvu4JS28WxI0O38t637xVeeJZ8Y/taAblPwddPzxQ1fmZeiCvtKQ
tmnkZy/3/UQq1nhgK5YcHblkdjDUv+CFG74q606cgG2GnsC660hiFmltvPlWWwp0YaYAhczQEjDE
f3T1v7moeFYlJTBsP/LFCUPGQFf3jGC3n0gtCNhdfBit2PvI66Q3dxCdrZaErfPDbo1+Vk9OC8DM
XmFoZJd9rOud6MywWBKJ0gEWwvjhD3yR9Jhzlg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6CCDN/g17uDgPb5uo/DyapeM7I4Cp++bTWpLwPsSWCozr67e3UVLUavvHI3XcCG/tkOmIza7cG4i
AqT1jvxWSno83Z5sIPqtMbKK+tia902lvGaJIR8BUYFwl2x89Pi+ZJubkXiuNgUzWbenysw9VIKQ
Gajcn5o3NDn2hpfcKAroPd/k/F7xwyd4LAvW8IIALz4NiCVoCAJkW22PZxuvwyAbqnSrSf4egCEx
pKV9CYDbEUYmHuezqE8VC3h15WcSGUITwdoXGxrXXJKm1+fEIWnv4THkaSczknggPRvnga+T3H4C
iwjfazrLLqgUxoj79hj5xz6q+sDR1e41lvXoLML4jTGGL7EMAcbebhBGe5q8uKNonFiY8IegJgPB
q/kchuhcQeYWDQ+HF6Y5FabYKK9IQGVRZ12/gm4KxhoJJWuREDMMAu7wIwsRaMxK9PJgWPM9f/Ez
A1kAZkdFDOk0FzC1TF5+CH9ZK04L3DqJdXDqBrr/zoPRVu9FlbPiO52TLn2scfhBX2rEH7s5ssnl
/Fat6q6bzK5hKZccag7MQd8AX/gDF1cW41DEQAKbuxLZlYDzD88/A+zD/cxAmfz2Ajsyxp21aKcn
U2g03nkBw03nZK0vUfdip3Qf7f/EExPLipmPh+hI25gi73BckED1ViCxwelKTg8J/iGvAzvOE385
c3A+PAfadotuPFgBrwctrE5Wh84mSWnY0E2EIyFZppvC5HCTkdZwQsh0kLTRXDDs1gIBW+w+7LiK
baD06lWQKkM+CeLHtU6gfImrSXK337juZg1mrNYXBA42igGBUTOtZMdXQWkk7UboeibG1DNMv6Rl
m/wzOwyQ93/S6ttYfSi7cG7gzNtx4uVxek8lfUmFTc6yVvMOg92NGBQ51dRbdJn9Zw9CbPy5Coeu
F8DeNv0gMabVI9r1LIO1v17vaIKO9tL0aYhLb/5rMW4E5VIJFnoDK45v5aFzf34GxMklOkMb3PVL
UvBNulit3jcHJaLUQhnmhm0A4CK7lKX783w31VADG1ueJY2vAhXTdvA7iVkBiASyTW7PifCgKLou
IotE4eaz/U4IYRLEgDXNBvJ+jbos0l8lf9BwjeTPqqMuGZjUsgUBlOL+pvAgC2spBAyHxrD3OGC/
rMVstBj4h+Dja1CBpBi4Of8j0+Xnqq73ZNTysHwAhuzjw1MLnGEOIRl7QB9bSU50jC/O98dTD42G
61gu4Cvxn8FhpGMEM8ivQsADelH8zSwffiFt9LzUc2nT9NSnHAX3ZxSHQL4T/QtWShZ9N1pisk0k
0vmqvdVf0NKcHpe6E27g9hy4+YLQhw4FI4CcW0lzOUSLm5HESPYqCDlAyxKe/Lq3V/r+AHAn25px
a9Ov1KzPUja0A0SJnpIWGt0UJ4PB1VVwLGe9CnvIRq/A7EV9icMQIAXXZL2zBGBURc/i+mV63zwz
FotfZBLVDIwW4vCnPTmLLB1q8Q2xwVUSITdD3kka+RmEjPs71lVd39yIwGUJ1MeskgWt96PN+qH+
V4l3Jq4FgpDka1Xphsix3/uKkU1YT2bLWOTivZxUhdr092jS+m1FtRmbJhjBNyys6Q3y8BLRVVy2
+/LUSa396f/4IBJHWTdF7E7slpOlZjONqTu9NpC/u04kYT7+iJg/ph7dZLjx+v9WoTOrZTLN93pv
iUZnIaD4fgnsjmo0KPXUhcfCiomshwjPCnopu9ZDoxPv9KAV7PCxjZQimwmbEMmcNgoGvHGqCqt1
LqAuqwWTCDevnbAjuXBnvqh61vbQpLhgdJPzbrY/Yidc+CSxgps6jWOIa8PtZYn0ccgre4Xe4kDG
ybTTel26mpr4CwTfkGMipW8UGvRRUa/xnDec9YsWmAjNNgg7/WMxyUeH7+pFX511L1R2lp61jMZM
GUGktXLTuyfl+IOs6VRAyw3B2TmW/bsa46t2okHc1HACyqtBGE/9CfQEbOxX8QjOTsT5ryAe2yH9
az4llh2F/Ndf4wbeJdL5YafbIQzMKHwQ4/8VCMT8FRlBKSB7kxsp93CtlLtitI1LnCsludV0R+6H
0k3RVeEpaTYe1iyd0MvhZqsvE13DDVF3gXSY87zjzWFBiCrIZX5L6K3DMnUQjb6GN0rWhfQtqpE3
KtzQ6BSjlPRD8TkE9JAzFHadjdRImOKF9waVauPf27T81+9ItDzehS7uJLhX+1lptJAZWxDVQB5s
qBh/E6OsYCv9jNTdiovvV4p7Wp8jZzEln4fMVbKCexdfDZwLwZ5XuZLJfw9Y3h6nzVr+5sxKrMtD
Vl9p3Cfr0yf1iix/0jbLQl+egB1AaHbXZKKMWkPiSZYllV9gSXPDxFKmB6pkgikr1ywIYgGQZRf8
cAeiSjatW0QD1yeb5esUo9NxW+niLuDwV7USSKAL4mo343FEcYaQVKxaFCJRikqsQr1cqrJrICs5
sRWaSflSC2vMclId0BD+H7wFmwASKbUKgmttyuiSjinaGO/O6/R0BCV5NFyuJVxQDlYFduHGqpQb
llauvUMHSZrF28X7wXFZ1oflJq4StEuQB5snL2Bc4mtD/YuYbD5Q8hApPP1hqzWTtn1Vyqjb96dp
dIQ3HUjv+UlT9GDgAekrDO43UFMpA2/KQh9Fbtosz8q0ZBUF7U9iV9mEZvZg/e/7vfj/qmQUcViT
qDHp5QhpmmGpxQN4FCo1oNXMd1/SPu+EJO7wT1yl8EWSNDVg4Bj//kbNzIIz9WqJC3Xp2SXDzia6
XX7xx6cTarcwSNkHPTA3RsuZ/wX5M8kYC3JgtLmcpMDDc8MW+c938PfW4P7NagMPtkHzusyom2RP
i2o2Y70A+adfyJJkQJnAWgf4hfRWKQ5LfwR8lBOwJJWPebst7oPgVvgxj7WEAPKcAjNP/GEXELSQ
+fOC3GhMt6s/6IKRopZhkDxwd+yES7l82uc+74vmDR3T+EmYb9hpDhHoBkYugUbmX67n7Yz/pVTd
ujTOBL1KZSTS6E3pOaX9W7TeqERF3JEzclR9oTwYKNMglTJINZLfGOVxHSNmLE+Y8rH4vmq3Lqmi
XOkGAuemMCd5HDuMgug1hyydEoNXzANl9ooluLTZigEsmhv0ZF4rDPXcGFX5C4Q2RhpbJGmEmRl9
JxIZHjBqSbBlIzj/00Sur+X9UOSd+Wk6eqDjVsuU5c+QswjkkdQIfPdlG+MUQtxyiEZ7cE69ad37
3kJuGKC7Irttntcw1xQrdaTyowISIJsfQIIVfrDOMGJc+w8Iy0WZ5k+86SJ/Sk8U8vH88m+3/EOj
S0XyX0MAwpM1uNJfwFsD5JJ91wyYZo1Xq4T/9IBPXoUkVjmwZ9E5Rimnz8RVMM0Cj+G3eifTW2uO
2WzIGrTy5j5V9evRqVitR1nA5xUMUfwKpjigfAPeb4iQFp6RHuerKN02p7am/iLhItdQEgvbA48n
A+Z2DZZbR5Ohm6CmZd+bpfqCOOm0LmPXwdvH81FTIDax8/u7udG4rg3DamcekUS1KpUFh7bG9J9p
JDYOsHJS+PGBaZE4n2SyW3AnA4I9z72mUOdf6rg1LwIEYpG9WbMYzgBDXkRnbfleyyXiJPamHlZc
P1eum/yWhb923jA5+eiARVJdxkEfqboB9u8fsMbMTft7Mr4lZgLgVqkg53I5QHDvjzPq6sFNI6Ds
QWSn8ZATqgphOGTwcegH7Maz4ptal8Fomf9nMRhP3WzAYGEH9lv2AVTUtxpu+nfGJiyLBNOj7cvU
VyXsjGrLBJFn5CTMoo6wMQqBKYpq/lt6c3cFh6j8KNN0Qzrj1jiOdU1DvAwANiLVQBi0+lIXuTl/
4hYWKMDU+RDYhsG4XMX2BXKAh9emLHm+HFteD41OiPJarjKptnZ/SkxVl3885JKcn4cnsZXCrSnX
JbyfjTXz9eFtGunWTwGbFXfcgQlxP7nmROMgrp8V5iSVuPb/X00Ae3enybaW5aVQUlaJ0gzJxeb3
LwgFsCdAR4lSsU5ljCL+UH7TipCQ/TE3YXJ5UsA5iYwa418OURonIWxVsc74Xy0oSg0GZohKkyvr
Gm7a5quGGxIVhWSK4EDRJW9tC7jOkWyWH+6VTwrNIFEFdX6dWzOkg6WDK1aqKGDzDzaPyPCyxtNo
rCArj/EVnpMmrSxUNCtUAnR2XMMIyzSZ7m3s1BdvLyUGfsyyx1shhyMlZ56AgPrNRetYwhanIria
YSnIGEF6QkA6lNA/mrBOOL7UCqrSagBYmpVjcHv9ibZjcczTgM1PBuy+lwqI7wjKbPZINt8G9C6z
Wbji/IfvylkFbuqIfpEB5/uvZO9B25PfvLYLvnOsRQqyHCkNk2G0OUik/DniCt1BdFv/jvUdQcY+
eHeZGCdMMBrPftk9c+0oD3zePiLQ7UVFB0yWfF9Eg2I5n3r3UzqirngCnSVkEhmh7JnMCjl0nYy2
mQQH6z4tFTu3ds2YRLoV0gGZncS6M5hdjHHfm3PATGxkkfdMfD5VAs92168+8VffT1PUKa5RVjhK
TDkODYfiMBD1cBVJbDSH3tRU9uzdzUDWBVkdPZZCdsqgt1wIsxt2YQE0iTdYNLm3Me+ILO1Qm4EI
3v2VW9FBCZUFeDcLSWSc+GSkSJ2q/iaWJQ1cyl8YgNN7pbU75FyrdevTi3qvh7yhMdKaaTr786bn
FifSjAUPUZHK7NBVY5NE3KBuY0ZBXf5ldHD8Z740lXR8jSPBCa+1hQHMD8h6Om2FGeSt08XuLToQ
RPT1Z7q6cZGOTk35Ij5IQJCCyXmyrkOsbr2Zj71viRRL3yMnqCuEZ0zXUrXDduJGvJEnuETOdsFW
gBwpzv19MEJDl4aKZLXPxlpaL736Rr2MYat3ayrtshk7CgkZMzwszrMoKJjWnEqG/cHgfOybUtFL
AWI3auSpIK7zNwoLrIjOSmzgAo7eo6rkbPUu/rmR+x7EtJj0SHlYs8pKe1KWFZO4IPCOpXts1baO
gMguNhDZvCAkkCuc0SYpjMoJq4Ln43dhIlMPcAL3bqgBbsqpP5Dtwitjc9AWzfn6DeQliQXBjLIA
l1fGXiwd1AHZT1zKec04SUZMYQZMrV5dWGR34rqUCbSQCIA5e7L/B8dPvwkcHIBK6Ul2G9IhqFjh
JY8OWrU9pFEC11iebfVQIqm1MBzE3hJdttjwx1mJvao6A1GPnzZtvVf/9ydOH6seMQD1M9f1YMVg
gG3PXAGb8i1DkMT4XxGqPGoa520vhVZui2+qe6rxN2wv2z2E6rco/pLvnbWMJQ2G6nsYqcQu9jPb
sdQNtyezkFQL+WO8M49bgFhiy3IBSvzNRpaoVaASBC4khcuMBAcFyU2mPQM1MqhtrdnGFIbPtQCk
IvhIQQWJ5joNEaRmH8vwSNbkjkEv7KTzrTCElK0TE7zssu/IELNTMQ1n/54GZ37wZdUW5OpX3Zzk
cvhxrkLgk6WOkZISM//zLLWZ2ynVx/AEim9SyHZnNtmbiyVneLkkbr7HocqBx9LoA8mHA1iStBo2
+mFU7rZo5qcGAW0HM7kdGNkEFkSfostX9JGcJZD4QOeVyrp1FN7RZnyBN6Tr3XZ6JhxwZNM2c1fF
W6URzH1zcV/Jcjl7uRPJsxGJyNVz8ex9tY+0Pwu/XodMd5h+ZEq+ovvK/W+oWonJ3PFzulKE0JMZ
C8wiG8x4o96TqJy+VZ/dFrJ7Kje/ol3p8ViofqsyjHk5gfJlQhG72EL0HVY+dM2pIEUgyQQC9iGg
eN56bWLlNkR5cx3b7cDGm8ijU+k+9npUpNh82YlDwz+laSUgwfH2ZnnwD+reNfmJ+WYeAQ2nu38e
7L/TU3Bj91IeGNHV4iitwh1hxqYKQznI1BymY7Ffk7xYtw+KsKt4Tb38E8xE3G4kHEEPdyKKlUJ4
URY5H+rTwFW2w57CIEI24YAbfkcoxiR6IG+Rcegt1Me+B8JFaTmLQXgCf2dOfMG0dtad6Xb5aQ1+
utTj+i04G/AVQNkXLpOO+RsJyQhwhR/wazqzJ+lU19HatblOXI2IJyItbvqnAp5hiEZ6QiOdKHPv
xmznzBr0AdCtPNRbwBkDRGZSU0VvyLOe4ihzXhmqBR1E5vyOlhS6NbgWcksFkmiyViLO6N0Y40P7
4OwD0ZLEmT4IgUPGQrig+TqAA/KtLF+JJ/YNEPBLTVFzuZvjVtlapX4kXtnaLBnasF3V4HML9S7O
aTAcMXsHXGlnJoSzjgAzZ45qbB95Du8HV16r1wfuJHCuVMOHx8FcP4dMqfsNDpqvDZi5N3qmYM/j
Kjer9mn+cn3/bH9NI2r76HvbWTb+oFoQ/taT1nrKwxVdJMJWgzCTPLMJUhy1Zmai5v2bWBR6BrrJ
wIludhRFq7ecaQ+bzMuyKVimC3TmZcn72QsP5TEZvNBgI2sZ+kvqS8Dd0gFc703OyuY80nALbtNG
vKIrlalbD/ASGi292tIHQBHomP3xtCH2AuCLVzu7zl4L2xl+yJDZBjZzdTPjIYiSyUl/ryGbdd1I
ERWYccTD/wChZePC2hHAKXNDlzLT03bnDPBbpZBNQkd6+d6peD0ZTWqCMG7/13sQzFwSMLSWpXJR
FA3M8QLKYvMqrePhsLntUZ2tekSs8otW5oD31/4sKWoFlGGa0/SBvuEwRK2LT3LiFHNZ7jLdBI4C
BerFxnCwXqdm05VaKZyVVNDmpTJPy8Tt0RlLSycxUdQUru4LtEk0DEs5O0hiebyuTYSDgmmAVc/s
zGQIFapRJo91A/seh16TsCCKSFuinD+7A40Cz1W9Gq53WtKdR+RjjBx14ls4Hz664yxArkwlzAt6
RTwza2x/SrPLd2R3IazkZBOodWTcbqCSTmTc96pcO1o5CD8wCbtPw8qCmUxvbizmoYx1V8SXFw6m
zAjvwLL2Sk0VNjMFvGLawn41mGjtGjHqmVfsOyPwW0uYUUISDhlI6P2ZWzgmJLkCNAQui96kRmkE
gCONpbfbM7ywcq9bb4lSPBZzKHnAd5oUNHb9Ip1p1+3CL5XCNMOojkrzE14Z/j+ach63SjekjBxD
nPAJd2qCFDLjZWH0rqdDmIY4+p2tvD/PAixBTBi4UOYlJU6qZoc5t/OjEWc7djML4RYusxkXvttN
eNmenISFCaHvO6TFCW4+/deTU32SWw4MXSl2OBUfSyjTOWvqL/vvfK8wHs5fvCXvqrBzyJ7rcA6F
OsQT4/qv/jOaHN5E8LWSBW+oW0GD+tA/k2ElFGjyUiWVXznGB9xHJDn7LxYXqB+zN3kiog5TJYKk
ROklV2K59hjH9UITi4HYwnimLdzWU1ay1x8WHvs61C7J8mYvPbNZs30DfE+GDqMknnIhLZQpyHnM
5HHJiqvv/S42z1RZU/TkPZFgN/9r4xlKNf4JSojRQ2w6AWyhy/vyFm13cHeAmaLhqkwKe8mh1Rbz
ngQ+ISHAfdGUE16TtXDeLRGEiTPAkMixgCqFcVWcCtZ0rJdHKTf+msGVvS+m6gfOh9L0Y6ke//bY
suBfYxVVqertgIq7jTDI8B0z3cap228vCeDMKXdlJP+izObwZr1e3S4FDg8HFgEqSUC1b0oU04E7
NWqNKkRHMm/8GDY2ggzuLTUEmsHwcLx8yvz0NePPTMLlvow6iKwelu68lVoeMXHoayy26RbI53QB
AtTqnJKsBz1guMdQj8v/Zow2tAkEgNCJQGJ8fiXRW+2BnRnkXoRVZpsfitSsPKFbp8UO2z6wiwGQ
NuSWLo0igcbK97wfmL+mCIIxiPSeiP2fhkC8FFS0E6v5jPmDFzEweBAOgDjLeZ0Wl0D9JCoj+1s3
u6zWUSo6X0QPCVrHrSfGTgZLo47dbSS/cIOX3eppXpuBsLoNVCM59YLBdoxM9CaoOaJQEoJssfqy
QwybOFA6s8B6+63mltMuJNNXaPDkE9P6L5xcwlziXKdkeA41iCHLRf0JAjsi7OmC6DpsRkLfrayr
4cG+RUDpxeRS0JK0lB5BL2oh8QYq2hnIWb2CX2zcM9ieCVrgKa60C5+ttDDlNF2KTAoCQnB9e0WN
zCW8NSmnquKTm6i5rg6p5v73hSXMXG4TW6bJEFAorGHa7Kv3N5250mAjwtD5FPw+OQJHq/K+CF/x
0HhD87UqdjJL0pXECM4z6Iwwh1jwb2t/lZxLzEdWX/NscTcN70JpZga1R/Mjpi/idGJFxAk+cbzi
tuQ6LNV1vkZmjZgn9XXwwzBRva8itTOyVRNfG7pV8bGxHSVNWC70sW+5dgu5OQevvbwXnKnwXMZb
nXkbAuhNCmasUHB9/cuvoZG/Ej9cVr2M8X0V2RB5R7/0/Y+8mUyZHBhVV7AFMgda/IZ8IuqtHI7k
I+54XNC/udYWviCSrXmGNK2pJB7tDIYKnO0mLpGHibDaVY24QkIUMxS0JQyveE9GeO5+JkXYjwg5
va2E7FQv8jFxrV9X+dPeD09U8HHJXkusmyQGrTxAuFw2A3HbisqbX2OGlwTSRG1Kg5lI/6TL/R76
oqhg6o07piSQE0XUOM5QmVmX9he7hGAxeGdn0gJd80HlL7FvbN3S+BMJFSun05eRe1g/KeMLXHKM
PSMQy7v4/tQ6v87QJdkPV69CnU9c+GaaUrFOWZYydk+4mV+kGuBFlP+c5GrnZpj2WB29BoNC+bBk
OqGsoplHBuqXJYkQLyb3HTwNQEbSbk74o7fPWq/SAboD7uPGiLMOFNYG0GcyLoLdv8lsgyGe81As
eXV17nd7t7cHhkV+cF2rZenX6rQTWUNeaiNMG4rFrT6eVCKRh018CAQo2zSEJedTiEAzqZfo+ygN
E4mjiNr9GNmXTPOi1UlsHeGZC0S1cu7u6symHtLELWvkzWFjZEzoAgt25JuK6kW4qE8qupR9vLgk
Ce8sujUA7w/RoV5uVEJcvhnKFbC9oB092mn9nOaV9ewnXgB6+A3hjFjPw+glW6HZFzxCiLrEiwnO
qqfPw4/nk6nwUILD+M/t3uUsISilQor2nMqkh/1uE4YkvV/aI+FpwjqHYiOgVuZFSTdPm2lVm7HG
q/L/x5+OBHEExk/hRE3FhzlUyg6m4TD7jj7I5srzjEtgfYuE2xzx7Xph57n1VVWwYPvJ0PpUmjpH
CsCGK5wt6cqMAQ8imb3RRTau8IJCTZNm05pg/BbpEZvhQ+ZoLSI7nCupXEy8wA2aDFqC7m8EOnSe
v0sgFdqoHM+E/q1STf4icO0IXit4qSqRWy7+OpL4gx3iLppj4HqGah6LU6dHQNaYUvsPWxNaRsOe
DY6pjjDBbxVCkhHBHDcEspqKLYflYJKIQVltnaZyAxV78d3zlCwESrqtbr2klcXrMppHlZaK1kDN
bxUjfxzvt2f3RpeMigD6cCvr7TqQR2r/fKEH6H43c2N+1clTWCoLore+JtyArDMTZN5DjSuPZrRA
RqafIMizKGSuH4yCbu9IK2Scuezv06oeyT9kjYqAWkZDzdXwSl0/OJIE5+pARWeIhM6INfvt0a8Z
D/Ade298oEfHfHSl7yk5d+vCh6Xa04KxfvG7SMEoH3PxbrTbViecodlAnPY4dohDnPw0GLCVTdH7
k8dx8iAIhhLBq1V1RFhfKqVQtlOT87T6S1aCLrIscl7mfUd1SvcmtBXe5FxFfO/Rwa4zGSJFRXwd
Y4K2UaiExETFPxAuySk5r0jmeBxkysEc6x78I2jotXskhwZZp3jWyoKJkT6cN3t/TzZWQlS8HdCG
BKGKHEqQ9s4NQS89AT3ji5zeiWRD99ADfsGQGl66jWrHmtvTEoj6f4/HqUcG72hWT5Qf5tEbj9eA
YADYlkd7tspZ6KjWV1N8QF5H1kjxj4XTzCX243ZSSTkL2iWOYhb86gtcc7RWpQHppFz/6sn8+nIJ
iPeqPgR9RDlcnwppnsF5F11MYipcru7nWgUGb+C9GXeJGRVCTbZ9CEUI0OUmawkzyI2KsHdCpWBs
o6RFDy9eCdVrPZJWycusNccl0KlHuHI+Kv//oNvG1rXpXA+jhBMM0nJtzfuDUPpSmU5spxPM0/Ay
Hcp1OflANDBgksTBSCQcmueqiz/Dngfhi1PatsaY74gLWkZf0OWbI6DBwMSmJe70wcTmdACXDEgJ
yZnygx4YiLXtSIkRcG30aYAJipsnukqwJZ8H0Ro9PQGI+EYy0OIgtDrTj4yVFYc2CIfHtrXpSdXf
qJFvejgxsFdIx2jaRIpoblwLVr+v7iFOz4sxVmYumHJQvNDHlqmou/8FBYw5pCGuX9d11LCWFHId
NfPthjDzyiCd0hNhbJly/TC0kZNZW7RKlQHScNE3ELhYwe4T2jgN5L/gvlW2PVWMb76ozP5biKK9
hXNlYrVzIcMJsFDD09lg8ZS+Ya3NqmFzlTxUDQ+n6DDOqyGJOtvRICdKbCnlogfstRJ2uKgf/csz
BYLJ5CA8mvFKMXMGygBzYzidJVZXtqZRxliGZAZCs+mYxmcSueHrOCdcSNqJJ6G75eWVZgcWzJHJ
EqjPJAIeTf3AD24E3gY33Z4HLu1KmcjoU1A1MpocTl/rZOB46BmnuXILQKPBsR4cj7HYtt1v6M14
WHNMEWFKeMQI+Cluvjgip0Xwk3J9KJ10fGkf+N2396OL2324L2cv6M9omzT6y77nk9JdUNvRErfN
Zz+S5N3M4PTKw18+MZKyAeA7R8C1PIJVv2g+xt027d7lvBrB1LQb/JsJYWcxPv2t5jkf+L0hBukc
mg0GQs/cmcj853+zusg2TUExgCLYt81ksnq6iCVm1hHj5ZtZ4/+rgvfaxZdZObH+CHvFuIeeLHiG
/RjneZMnGSsnTGHPyMA8TP4MFY5Hk9qO9NA4MMbOdefjtmHzA1FCpWOBEOvJZqsFHLHL7MGr7auI
UNjUf6x4Pnb9BOmIOqJ0WRuYfDhWp8vyEK22h33ZG6EoHqKe2dnaeBCixdEbMx6sqOdxbXuKLPIA
efAu6SDJk7DuYMnlUHpxS4y+hx2F/0oRlVGzheSwAYFhhYpSM1wQ4Uyq6cVu78fbnmVGpQWUU/QK
R0sB8eS37yMxyzybfxiNOLqELu2tbqTMVXWeQUFf996bdlGDYouv8lM9excqNJDvPwx7fJRcs4K2
Qv6WjRFZavHPZd8C7D6DM6bsQGhNBjubXG01xTZY4cb2LdIBHnK84utJNB2oriGk94vH9tkEaaCr
WmVrmtA6q3YXfAl2NQYtIeqt4HwQl9baPMEiwDgV+rhsJcoyrMxxcljhhh9sm2ZFzb9vU1WTKsnf
oXlw2W36xw9i3Oz9rw4OpvYzp6ep8M1bUJ5GfvidINNDFg23mG+Jwx1xc3eK4/jIu14gz/ebC+8r
Q6Mzt5nk6p5GutTKWMLD+jp93rRahDOfvA17VeeDQLM5CPvlzdWjfF7aJty9D+ymHFCgDiR55IRF
e9zpHqAgw4ofrWNYqL1xqARCPG0No7SDAm2afnl2ayCT1zdPCZ8DuBMc00XWjpDTEilQJt1yMPHY
u3/bzWM8HFH0NR6dhpgHzGA36CQDxsLykv17Gp7XsqMFNFo8mJPfmhYrBgsWUOr812Sw7h5Sw4Ja
8FT87jshLHEPUiGld5U7MeBrAUmyZvGAswabjYeXIVbB2xgOV2ipJsVf7K85pBs4WUgHvySh2G9B
jDJzePuda0LM1VsxWm9OjXX2ETS7Hq2e0Vhp7A51S3aVse8ykqdjeAD5x4FvET2u/bjhsOKTkv57
V5fh3aedYBELuD6VQ26W/Q6DjcWD6t6U47OmkhFQ/sq23w6Hf+JUEpXp/zRJtdD/C2NJPGm06QCQ
Mqxy9pFOb2W+F1XFxgA+EGv1/+Tr6QhJigdvP1JX7tY0nZQBZLnponaz2ODlDDND5VofjFxLdEN6
TNZGrkgapW5+WitqkGYTxT4BXtjB9ar9OKwhRV6yaZNWrVb1h1wkmN21FCBRKDlbPt4uKH6UiNPE
QqGg9q1/WAj4kWTNk+JZe8AqMGciBtITe3rVhy7ncFRO6tPTom+ggkL717/GDuCabNX4KxQRMGQK
F+UezyHLg6bPTz7G1JFWoN8jflQPZmB2e6xfOl6EJ4HYKCNApo5pAw65Iq6Exzj5s5IXI4J7tyoZ
uecWtYb5DcUbWwRphZeHiYH2PqGblXPD97cDKG797j68P1b/TVImZ5HyropSPi61ZpmPxSWgu9V4
YosLS7DBOMBtMJL7r2pamo5i6AXRQKx3DjO8koE0Y9M/3zYzHI2SKoonNbXmb/kgrPONfUTxv5tk
+gh6NVnIhJil/H6uuLkxuyCwBF2d6JSCIhC312WvNyOIiQTHTLqCZOGvdUjDzCpPKylMwEAjZnp/
I3h3PuYv3E88ANS4v4UpbHq3qMIQOrn91iAOngbASpUP0O82Tkfyarhngm9ii//MgrRax1GFqC7J
z5Veor7cV5eE/UvaTqP/NGS2Ofn0Jr97jzJ9f1kepGGw62XYA2MlIipDsArN/S/zve8iV88VfcXJ
fK+wxtQ0g0nIUXmTShKpvo5GAWIUm7aHM6409/F0s5aUo3hQCn3rY0TePvEYaU/QO45cQGa+/VUD
J36f5viuaNujxz9tedNO4SI5veZjKR4jXYD4T/kmtuUOEL+YUIGxogX4JvgKJhnq7Jd/yeXGAgZO
44SuymBSNV5zoNDIqEhHcvxlz4D422X0nw0JKLesANzD5c/b0libH9Crgmo4+sWlEbEHcMGNnlOp
DuNdYPymqWkK6Ipd/YTw8WBFWYjirjSOf1jQmPI8A/2UcSyZCK31yOaop33zsXuEXp1lomu14Dm2
SDDw61zVf7MDPHOoisMnE6ws69Tks4bRERtJsUuDwPnU+RD7T2oO+08Q5KZUByntIh37MwHHflkA
PbmE+sdTXsdYFm2/g3xBe+nmO81nz4uRQUejN6qW5JBK7TCQ86YGoA7jU37yi69NS9+kPNysHd80
UYK4mFVXFSyvGwKtyjlIUg6c9kzin+noIUpu/1gj7AeIuEngxt1hWQU+1VvGSywdBxN3fYDY9a6E
BfKtGdYeT+AftRJqRA/DJtP5vG2FQcCOrfLcDAudQ2HvnbAD5z4DQ73rpreE8tYvHsMLYqAxlTyq
8woLGnuHxmnB49g0fEUGxvkkVjF2HZxkFbqkC8nk3YqbWH9t7aDeQzoRpMP3uPsGdO3VH1JDsyZ1
+Vd+OzH0DGSkUZ1ASfoxiS1Szlp2YEHOIfvbHbl+LTewrvyf8EMayvdnfjqKsIflevjdCGGgNjjD
vaCmjrKlXoSbPlps6w75YgiTIhl9z10NAr0ImnPhEKKfivPxlMDt1Ia9/RCYmxyPFb+YAxHNK0kQ
NQ1IK4I955riuYsIsIJjL6C2VIL4len2skf+rgOZh4UEuHWnfQZAI23vr21bOMC9He14cpdYetpw
B3nY3lKqwwU307fek9VXZL3lwo2jSUt54NGfn1PRCjbBNPEZ0CnkXZupJokvHiL2Z56pRfBmqXcb
gGHbL3b1207WZCGwo4rzwcnMZS+dv9mdmh2/KYmLMqSv9ulA1ukdTmUiILNv9LudopPWvZuK3miU
QeGDtI1GSxr3guXMOfoXnekR8LZ6rQi1eu/8R8Aqjb05ypN+BVV2hj3NEwb21tbLHn83PASs+ydq
mbzwVc2sGLqQPji6bCfxaaz/DSkwIFPSAsorVbR8V+wM8df6K89rCLGOvqbzovV84J+/dydya3qn
p7w7jBsuwFcdTCCo5ze6SONDWB1mnJgB2Rxv5ns/PrbEDn83mv4VFa7J/KzIjN2MgBfKiaqu3Nbb
45kQW0k8tBMa8OsKQKVTSx2hyojanB0kTWQjvbqLo5V8L79eNwvtUdcRSKMUtHWmH69t8RzS57U6
lmx42VB9QlrlmcKIDnFHnPJGxHtI1uKeBjwxH/HCSWWskAuowWYAdoBrcBgIyVCE9LxzXFgA2Ul9
nRu6VSSfkFwgfLCK61WkejKNOcnQHLOgFg2aYosuHI3d33NdImlErdgd8TOMO8byrKoWNMaUtUV2
zRNs86yoDU5FA+vvlY6NLtT7uUgUcbwSfCrH1gZQl6MuZ4N4pnmWs0d3qYUfuAHLA7bA/AkvgWKO
hOl4Q/1h1/eKLICczv1VA4nEvG0JE1BD2zEc3/frzPpHHiTx5/pKUUpWHAq79ZYtRwsXBC9+qT7a
pSsC/NwZdT3ZFmWFhkPlcXTyIyhUjFiih81Fs2zj/ALNxiLxMKEBsVQJd4ae21xrQxlaU0jOGv32
884CT7mChgDwzZIpAv4IVzNfRIGsKp8wVGdOiOnDuNmFpRwOTj69ev8MhzCuWQmxi0HxdrVt1WIn
PToABH8oz0eWGt5Mn1hcsOv+G2oT9n2rqXU2Dj5ES7ZVaRzVvQWbZ2yRvPQV3c8GqK+BjUWUpmJR
yRkQ+nUSz9p++vMoOPT9Wtl9ZMTvgTbFnc6R7TjkRVl79MUlFD8Zj37BptdhAG7ZT2FZSUL8OYIa
coy/DVe4idACbVO4z2/PUoqRxM0qd5/QUiDu9hCuokYQsuxEJDLx50U1WOpEAId1y60YMj8tRipU
hQrEMlWvSE61cVQBJXispxuwTYvvps5EFeT0fGcZfMvsyEkaagScYtpPBxuCRYNRAosGh9YeWa1X
K4FG3a8oePjWk3TJ84V4j2fIzd96er5lnhI17nkvo01ZJeDksRk6Gdq+LNh2JIuXHN449wdG/8BN
6ROyXtIS0ONO7eXOy+ONPIRJFnfo2OnvcMNnmrMrvCTZOboOzT+F0WzAzuFzNyMLDpu+iiGYGnVq
5B2w5tmRMq5NhOxtjGL7MzAuUnMWIKA0l4Sx+UfqYaOth80YORb58+TKs2XXMss7UmJf/aNzn8Vl
tQ0iy7tdiesrlehvkR3V8R/Fl1qB98gnlq0B8VnSZq8QGh0HPb+W6FJHEEvRkL80WZgc6D8a4W3I
q94KbMOw4cVbe9uOw502AxkcVyd0QRfkbHpaYufQJwGuS2WwgX8uXZjVhLh7MlW5fZQkhjyK1eEM
RKgtpTAs0gCnnxRvSEH0bQNPDTmNvYvfg477WSfRAqBbc+V+LytMKUCxlZivaZ2CHuSDAc4Bp0pi
w0LV6hOXBmejR3D3atRmCs/9KgZHwWkEWW7ikRcuEIyKZLldtlWidl8EUAkn8YpNVHf3yhUr/rvh
tCPhhUaFTDlHrw4VTRkbko911IViisQM7+e9vJe4HbF8DIFZmWqesQyfv6qiQG/adSj6U4L+fDcl
ZdQcMPwKiB84S79oUc650RFG4hFnZghiKrW5EQ2pJbNTr5tHUqDXBA94sQx52QIv5daWC5c/RFi/
xws8k1Tl0ujFgZTpAKVWR8F9EoUCPqWhVNDcEsF8TF716lv5zcW8eCNGXcoEL7vkDpPfYWVPtIKe
IAzw96o63oGj3jiQ/dxK0YtbNdpWPe/5edjGz/jj/Bs3ZU3eaIQBkL2WZW1ypuqKj7l/KPND2lBF
t1eY4BYgj/rUO/WBOPSO4t0NoR6N+eLXawcHmbVICj8woeM0mC4JIXLjWuISyFkLGqvq91ajZC2i
aylzLKa/tT2JVdgt48hsN2PV3s42yqcx+fYr8/Ozz7neXEHF+yGXxvkwn2tvoi02aS5+0rH0fgyc
oclwSFjSYYBEmgDKvEeZ34O9c0RLPzP8EphB7wYJOjKXizf7HOsi4zQ5rduyjMhJq8jvHHyeW0xV
5yE8CbzzbB0zhRTCvzrwgBPRxchUaZecF4dpm2NBXsh8LeHBSuoULW79Z/xE+8YUEWe276aaP7/+
/L1757Fkj1tVp191iRcL9poYpU0p9RHhjyfD9DrZTAkSxGIOGuOXZtXuKbrhGQTFayrnncAJ2Vmd
tDvrElQY6ULWC4QeIacoT2oB4pzlHP4tDWQkZDTJWAcBsU91+yi/ccn/DsfkwyaF/0h6KrJNP6tT
b5EjmLK+8vwAlujDZfCeP72xl3mBTsvlHhXANrE3TG3rAH0rxZAtTQufxkQxlyzdPmjvQQmGtFZt
Bpdi4YIvPyie8T+291SmIU5wTqrxITgZleYuQWhwojPN5vXugcOwqvULRwxuaSvqgMhURcDNdYfj
ijBFVh+a+TPQAhQEfwZBsuN/nGhKb2GFKiZnT2dTTU6/acn989sxr3sr0qT1YQ8JmQx8WfjGZ5ZQ
3a6KEwPgnXKgmv5TcKIMuzjg76vDfHOK/JaHNIoJY+0C0pyd0b1LdnfDCQss1BorINmLjPrLo+uW
UKIEvGygRfi4tLXYRWxhmqDBK/cgIEZWcWf433bRnXX7OT/k6rsG26ExKAgo3uVUUiSMYVKUSIOi
QwobCYLFOFeItaVrS3Q9oEndvmpfrM9g0RDQzfmmMm47HTLbmlZCxthrwXLjn5swUQgY3ohVd9Uw
n449mdEjQuPKVKES77ngBQoXnwdSJuaaVXzxxZtWD44662uOP2dmIrwlQ6tK2IRcwCAth5r2GAng
E1A4TokVwYTeWCP28KCasdpapXeS2uixeUBe08ySnHFX/AxNGigVFZRMd5mCquvXXoVHKn+XOHp0
Iy92GNjScddtwb09ZBhvfIF+MqmwBjYn6FTjtKrsB5jwT6D0UrzsZSw+TO+dDRcO8e+MjO5vIKN+
XMDsxaHcLdyLwmch8/8kFOOSVAYpRKpEzvWdgyOtxEqAaN0w397SsyjjTRsLNxe8KqwZKT1R7gF4
vCSuNCEtSF7zMCa6m25UDjahdNEYszsRx7KUmqKnPj3390hpq4teg240gVqk115ErTDdehnIfsv0
zyAgw3JdoTesSI1DrGslseNwvQC0Wf3EXd3MJYrozarHVP963+HUihb/+5EPIGcMFssmVAku+eQo
YR9CmGx1a7c8r6dM4WAG7zDYoR/990E6Mc2vF1thNo3wwmyofyFdfWsLcLS9Xe6HzhBS8mgzMgb2
RsYsY1kY6g5gfbikJFOBdfe1hIqzPTKG9fiM5iBDQ6zx4+eWBie2ykfxPnj3Lu0PqstRvIs8e48L
G4+/QF7xiMFzEnXSSlTTWHElJ4D3LoWGHNLT+lycjf2Wy/S5/uHnTQgguog2V0vxa4qM2DY4tZWJ
06KcSwJa9ZdvXQ32345BUL43/hO0RmEFT7XEpL2n5bd8r6TUFkgQl8N+4NORzD+jOcvFgXjeOGX5
uccwrtcVZaQBnwQe6J9ADeSmvvC8cqasKn9ca+FCdqYzfb6isqfqvcfXCujldXjdfqW2Kga1qy+L
6cX8sipqMsqJzRkBqhRVI7Ib9Pqt/ZQ6713xIRGbpjpJ/nwGTvfiB7iB+ExwDfsW8GUJl80eJJQO
U7m2uFPnTTfy9GSse+/ZNoYz2a8BNvbYHZZKMnhB/f/QT2A2qYLvUfOUwK2vyr8zvQPC+qo4uw6v
GlfvLrGz667ufqdJkea8j5PorjMcnpZ6L95fTG491Ns4PwEstwPbrU6EkXcEKCsp2l9Y4pj4IJ6I
mt8awuhT7o9hjbmL/7npy8u1oC3z+eJEntuOFcXCauhCJzWQyIwaQR/a+LIvrGwX2yYT56Q0A2Oy
blQGWXSvNXI4sUr8lnmt4FX0xmrnFOiBQXbotngR3udJNvw1jBFcPIwEs5nowT8fvfFPyfHt4nz4
U/Tvob1MH+nGqUebD3G20zeXbNLqIcxZ5jijXk+mhK/p0T5/8PZsJsaX6QWwNaFG8Rv770tkMaBY
yKxhgdwRz415BsAOKnLdInSIt5rOdhpzTfCCRRwL7a9xFdfrwe3yGGIUh/YpMCoiDnxSPOXDf/Oz
88tcA5IZXRLT/qbxuHTSfQJWBbU66IwWPPk6GPyivPNf3bWh/9iCauz0t++nrzILDUQkPhaLsZOO
tvwYCCTuhHMNdfbjy5uERKjizP0fzERpzhBGv6pIljf2AkamH6MkUQ+5n+zIEannqIt9mfLSle6g
WM3fHfH0QBN2nDew1R9h2YNbZyIwiXXUZrfKqwtiEk2WXYEt60dO5wWhn6l/4Nug1eMXRYf/m1A4
k/khhxnyhqerDXDPhkcolKuVWMFu7+gTCMAH2AjaLyz55yDS7Izq5/HqKgLcZv9jJno4k+xNYso6
/M/SsUWw+FHJFXI4Y/22gLErrwUO8tKrueyyYwNll0wmn/x/Ch71e35tgAkN/L/2p30dgXwrKUJf
vlViZ4xmnqE7d5oF7OUY7W9fWOWu3zwa0QgQD5gCN8c4nOeKBtt4G+FAGur+9cjjh69zNbJURXRy
ZoJXOwS2cdU4/9xIsdr8//8VxiQU3FFAIqV9s508v7ez2VciNaRbP68+R9uTugteR2oa32ElqdSZ
olauk+mU+D7qG3oilN07recLALXyZLiMB6Are49SnCJlE93AwLW+6di59fWQBzwGHPpgTHpXjkX4
3LVjWtsXA7nVdRz16hGbep+4etwOM4kPtAo/eFscw7WuBpb9++Fe/XJMF0NJwxU0u2/3TGgpgOtO
dCXmrsRv+mI7+yAnt7BbU/GZnQkjNXvZejxcFRVq1Jchf+zEkrsBhzQVNQbfzpfD2R5fa7ZMOV6E
AaDGwsCcOVN1947RgWQVd041ZfBoCHF+KuYSDXCKmmi+gBlXRu4E4AKPlJ03BPpFwCax0gSSzLUu
6tyqBwFt8elGFJzxILjFl5DVB+GTBT+i9uclwtMPmQaIYvT4Etxn+D628a7if0d5781UCMHF9U4f
ftNtB1Ja6ljYUyGS1PyxoasAyDOEx3fuJHFBF0EPpDESCPBu10JZFxFMMzNyddhSXdeB3h3IzgO6
VANBIgaAmPd5lELFmFuFa3pPo7oavt6CQAdPOyOd3kTflViFnzcvYOeBBkbAyDTPaSYNA1uLmTYW
FRh1i6U2LRkPuJS1ZxSgrhp7zoHeyIv3TPtinGSUopMm7/FEsn4pygXKHP90Uj2jEzDpQqCs0z93
+s5o9W6Af2Gzy7exxEDLpp9anEdQsRs694eJASH9Ct7zQQgdOTcccD82RajGQRugUtVeFWmreakf
q34IuzgPQzg3jQJLKAty08TFmovgyI+Tx00q1LsKSHNO73KGmLhS0H7iScq7dNYENiJUsQSgmmBx
kNCP+36E64gTKwyLV+4AgYqNLmmEaVK1/mLKdWT/IVLmeSBpXiO9BA+KJNeBIRO8c8HCn3B5YX3G
RV/kLS8yV7ZMXYE91CCaJx/02wQZQhG0VGzMN96f2jLNeGgLSpXDLOgPK74EKT34cPXI2nugBBhb
oR6G1iDmT2B4Ns520SF5kxwHGCv7rtQDeB4vpnGUGJ7p0E94U6DpvsFtBNzUVvnuE6kLqQ+SaA71
/z8OZ/PX/+adQj+HLB2Q4qE2yNQU3w99NyjDSFb+aedE2MwLJyXFCHUn+EmrQyPGg/i+ZtC6bDt3
iIZxbPzFYddqTG1xw9urC1Mah4VyzMKuW3sAldoBG4g1mqQ/58LhHamOHJDJJDkFpFpCPuTN/zfO
k9S37rfX9n5spMT3JO98LBImioX6f+BAvN1oI690kdTK6GTXBJZWAHmTd2HKg84zUolDFkYOlbyg
TtuHwV1kWfkvJHJ88HWJGq1EU6N/rltACwPDn8S7ljwSP//Hd14SCi+L6qt0gziAq/PVj2E9zsv9
dKYBzDjM+pGjkgyJs9j2NRnFcCbvu09A1O16PH6F8JPLCWBRtViIbAyR5/K+25VqHHwqsnolfjVL
lZNr1+HD+sPjVlPbUMzffU47/VCEmQvooLOg9mMuzy2F39PYX7zFsKRuhLzAeBn6nLwLpC02uNWC
UV2Abk6H2vkNMkXMDd+PGpRvym+NiWMKUEPGPbX6qLoZTxc5ihDNiqC+q0DQHsjWso3iggtP1p0y
6vcCgJHE4whtmOdl+H7VF4yT/HonaCBp5P9jzsqHCeLDqq3bqLn+RrfL0N6C6Dgjp0eauQeIG4ON
Y+3MAz+ji06Z/RUO1GaRWAoEIJepkg1chpg1x06gNRiUsDRUOxIf//qQkXo3XWafYoBCLcMLlPUn
Kiyapub48tmFubntCmfllDYALg8HlEUMOkyBmWIlNd7wdKiu6/xLARQPnH7N2VnIAumDVl7hDG3c
sSpmGMh5mQ8l4QKtuuYhMsFJJuhmSMsU2cKyps3Hv4PqylJBPut4aJFOgKDJDFFritGazWQP3bq3
iiVVPDfkLGrCJ0KreLuFCk+EwxYSASDxipwNUa5OJwFmDoCQM12JRpqPvWQQExRCc220iXdgDaPF
x+gZWnp3TQULk1lXEPdTluz7NyODoYzr4PvVitwxONrTum5f/YnFqBAy5iH2qK02f99CI2YO+kRy
3Hr/RSC0xrga8muTZfsZNSV4WsGXQy05BZxvE9bDP2aYZehTuj9Y4qlS8d2wSsfGfcp3rMwgeoB4
sAKIpCfNjLF+J/5yZqxyEHe6pGhKMer3VHzdT1dQgIFHaU0eRZQdomDimz9MB1rf8nuSy2BLJHEm
e6f7DU5k3oq3J2YkjrVRGcSC04dWr9LRA+XEZtJoXPivqGcWSwEdi2IjK8lE5gDNfVCEo9CtxI9L
IN0bpFrTPuswJegDJLno2GSPSSh4djWZ3DCf1S7XMAHA85MjcvcJO++JVuNqVh8waR5QJ73p+Fs0
UiKwXSXndljqVtJzRYpKNvlsV8Js1IwFMtc6rsLZ9xA0bm29mj5+05vtoL1stcz1/auf6IxB+PMm
3Qii7aMQTFhiwW9iA0Fbn5NsBY7Ddj8XXIdPulGkmoGpmp4J7bi5eH1BR3DdHl2NHgg1XycVoXp1
iloXXwgaZE+EDhZ/tYvRyHUUNkk5eMaREMR1U7zo4nnWkNE43gXV+KRlESjOPrCPSYnwmp/N3NGC
qDVyMkW6Vyqy6mG2JsmvFsiuszwrt4ZPWsxgu8lb3ihHynKF4bKsUNCnUzoPTy9Zg8XvxBJ0lv7l
FEv0nEu5JY6bqQTAdpwMLszkTq/KscOlV66cLgobP5kYaCrUZEboOtLPdQypociwrX/XDomclwWN
EmbuqUjoufjVvm+UGrL+9J+7GFtppfjmForO5+QTGZ6Ii0q6AWH7tB41SZPgl8QyatKtFb22MvBL
RoVc0Qk//eM6d11wEHtJF2cXqa2bsjw5HfQSGcC9yuiofeEvNSyW78eKoBfHXtEEKnjlrC8UCjs7
L1FCf6uLHqScxjjA2PtT5NunUsLoiArL+T9ZDYi0sn0QFNAUsPu5+H76AomxkaMFzNx5z4dqKjoD
LabDFcILut8AE4h7//8vxhqq1q1l4FjWzhmRqBzdboF2kqk641pfySsMZswTjWOzUxBOEnBIf0PF
t4/Kj21hTItijeIilEVeTJjMpmpyNIMK+C3TuJvVPUqabbYLHNvjH2cNTd77jjNTevjRtGQxbfQn
S4LY54Djkv1vT1nkC5cA6GcX+Y/w4gbYpmLciyHguhNP5Td+F4m1TkVndULEQ0rJsMD5St9t+Vyc
B+51LQNpy7rh5il3UTIff7AstpNwQwNihcNReMOu/gFUBH/Rkv0A/acQkVnzC6pR8tvfTmVRQW7E
Uall6CcxgbGy2Ezc1ylHiAJSIY+zyzoVJhzA8qMHY6d+u1suxILVs7wVmwOafhqR+bAlyKJR6Nor
g1k3t2flt7joLWkDOHse/vYwdl6dEL4ECA9eg/oZbFH4Zk85/QjOvKeLjYvziRQMnOYDw0PDxN1D
LwQhj4RA2Y8YL+5Be0Kz1pM6E7IRngqD/CwQMKVF7lx9n8gzBCeQYo01WQAVbkNpCSofHs982zqR
KnN5rfJTwzQgkvnMJAQ2a2rBBvev7QVAs9WkGhtWrZdvz8CAFRakYgkUDcz/2tTQ2Blr6vTiYH3F
1J0cFZGpk/DcxYoW2f6Fetd7OA8NyefJ9+FMg9J0hUlaoQjbtwAkv01d9MsHtexI4SnEXmC1tKnP
2YbmotHKd/Geyc2BQhGzuYqZZKCM9F/J/XVSyBmYRrLnRBj7y9J0m0/ojL56Jkhja8FJGOSMi58I
LEtBVkdkhVn9Jw2MPmmO7OXAWaGl4jRv6IcoLxHkU7jjjBNZhqNZi/I70uoIeH6ybldeNWA7swg9
JgCGb8sfggpcpa2lmG+AOWXOXNOI4QnR1kVag0P2oyxu9n8qhapV8j071O0tWz8fCyR6W+eIYUm8
wQOkbo+o/jcPaWN1OJUQjPUtDL0vUjGbf9FesEXEiuCGw56WClJqqCETynwxrcNilgATALV5PA8t
/MjYRlMW289tK5+jDUMLI/erCJ3gnS1BtkF/jY6r4R95oG7mjGZzxH6O6/a02zJ8lppWh5HBaIqZ
rLfBuCsFNr93uXe48Dq+vU6xDgdUrUSZhxH6hGns8hebKQD1Mg==
`pragma protect end_protected
